module anfsqrt_sqrt(query, result);
  input [31:0] query;
  output [15:0] result;
  wire [31:0] query;
  wire [15:0] result;
  wire [31:0] \eps[13] ;
  wire [31:0] \eps[9] ;
  wire [31:0] \eps[11] ;
  wire [31:0] \eps[10] ;
  wire [31:0] \eps[15] ;
  wire [31:0] \eps[12] ;
  wire [31:0] \eps[14] ;
  wire \genblk1[10].inst_SUB_UNS_OP_n_736 ,
       \genblk1[10].inst_SUB_UNS_OP_n_738 ,
       \genblk1[10].inst_SUB_UNS_OP_n_740 ,
       \genblk1[10].inst_SUB_UNS_OP_n_742 ,
       \genblk1[10].inst_SUB_UNS_OP_n_744 ,
       \genblk1[10].inst_SUB_UNS_OP_n_746 ,
       \genblk1[10].inst_SUB_UNS_OP_n_748 ,
       \genblk1[10].inst_SUB_UNS_OP_n_750 ;
  wire \genblk1[10].inst_SUB_UNS_OP_n_752 ,
       \genblk1[10].inst_SUB_UNS_OP_n_754 ,
       \genblk1[10].inst_SUB_UNS_OP_n_755 ,
       \genblk1[10].inst_SUB_UNS_OP_n_756 ,
       \genblk1[10].inst_SUB_UNS_OP_n_758 ,
       \genblk1[10].inst_SUB_UNS_OP_n_759 ,
       \genblk1[10].inst_SUB_UNS_OP_n_760 ,
       \genblk1[10].inst_SUB_UNS_OP_n_761 ;
  wire \genblk1[10].inst_SUB_UNS_OP_n_763 ,
       \genblk1[10].inst_SUB_UNS_OP_n_764 ,
       \genblk1[10].inst_SUB_UNS_OP_n_765 ,
       \genblk1[10].inst_SUB_UNS_OP_n_766 ,
       \genblk1[10].inst_SUB_UNS_OP_n_767 ,
       \genblk1[10].inst_SUB_UNS_OP_n_768 ,
       \genblk1[10].inst_SUB_UNS_OP_n_769 ,
       \genblk1[10].inst_SUB_UNS_OP_n_770 ;
  wire \genblk1[10].inst_SUB_UNS_OP_n_771 , \genblk1[10].inst_n_707 ,
       \genblk1[10].inst_n_708 , \genblk1[10].inst_n_709 ,
       \genblk1[10].inst_n_710 , \genblk1[10].inst_n_711 ,
       \genblk1[10].inst_n_712 , \genblk1[10].inst_n_713 ;
  wire \genblk1[10].inst_n_714 , \genblk1[10].inst_n_715 ,
       \genblk1[11].inst_SUB_UNS_OP_n_771 ,
       \genblk1[11].inst_SUB_UNS_OP_n_774 ,
       \genblk1[11].inst_SUB_UNS_OP_n_776 ,
       \genblk1[11].inst_SUB_UNS_OP_n_778 ,
       \genblk1[11].inst_SUB_UNS_OP_n_780 ,
       \genblk1[11].inst_SUB_UNS_OP_n_782 ;
  wire \genblk1[11].inst_SUB_UNS_OP_n_784 ,
       \genblk1[11].inst_SUB_UNS_OP_n_786 ,
       \genblk1[11].inst_SUB_UNS_OP_n_788 ,
       \genblk1[11].inst_SUB_UNS_OP_n_790 ,
       \genblk1[11].inst_SUB_UNS_OP_n_792 ,
       \genblk1[11].inst_SUB_UNS_OP_n_793 ,
       \genblk1[11].inst_SUB_UNS_OP_n_794 ,
       \genblk1[11].inst_SUB_UNS_OP_n_796 ;
  wire \genblk1[11].inst_SUB_UNS_OP_n_797 ,
       \genblk1[11].inst_SUB_UNS_OP_n_798 ,
       \genblk1[11].inst_SUB_UNS_OP_n_800 ,
       \genblk1[11].inst_SUB_UNS_OP_n_801 ,
       \genblk1[11].inst_SUB_UNS_OP_n_802 ,
       \genblk1[11].inst_SUB_UNS_OP_n_803 ,
       \genblk1[11].inst_SUB_UNS_OP_n_804 ,
       \genblk1[11].inst_SUB_UNS_OP_n_805 ;
  wire \genblk1[11].inst_SUB_UNS_OP_n_806 ,
       \genblk1[11].inst_SUB_UNS_OP_n_807 ,
       \genblk1[11].inst_SUB_UNS_OP_n_808 ,
       \genblk1[11].inst_SUB_UNS_OP_n_810 ,
       \genblk1[11].inst_SUB_UNS_OP_n_811 , \genblk1[11].inst_n_708 ,
       \genblk1[11].inst_n_709 , \genblk1[11].inst_n_710 ;
  wire \genblk1[11].inst_n_711 , \genblk1[11].inst_n_712 ,
       \genblk1[11].inst_n_713 , \genblk1[11].inst_n_714 ,
       \genblk1[11].inst_n_715 , \genblk1[11].inst_n_716 ,
       \genblk1[11].inst_n_717 , \genblk1[12].inst_SUB_UNS_OP_n_822 ;
  wire \genblk1[12].inst_SUB_UNS_OP_n_825 ,
       \genblk1[12].inst_SUB_UNS_OP_n_827 ,
       \genblk1[12].inst_SUB_UNS_OP_n_829 ,
       \genblk1[12].inst_SUB_UNS_OP_n_831 ,
       \genblk1[12].inst_SUB_UNS_OP_n_833 ,
       \genblk1[12].inst_SUB_UNS_OP_n_835 ,
       \genblk1[12].inst_SUB_UNS_OP_n_837 ,
       \genblk1[12].inst_SUB_UNS_OP_n_839 ;
  wire \genblk1[12].inst_SUB_UNS_OP_n_841 ,
       \genblk1[12].inst_SUB_UNS_OP_n_843 ,
       \genblk1[12].inst_SUB_UNS_OP_n_844 ,
       \genblk1[12].inst_SUB_UNS_OP_n_845 ,
       \genblk1[12].inst_SUB_UNS_OP_n_847 ,
       \genblk1[12].inst_SUB_UNS_OP_n_848 ,
       \genblk1[12].inst_SUB_UNS_OP_n_849 ,
       \genblk1[12].inst_SUB_UNS_OP_n_850 ;
  wire \genblk1[12].inst_SUB_UNS_OP_n_852 ,
       \genblk1[12].inst_SUB_UNS_OP_n_853 ,
       \genblk1[12].inst_SUB_UNS_OP_n_854 ,
       \genblk1[12].inst_SUB_UNS_OP_n_857 ,
       \genblk1[12].inst_SUB_UNS_OP_n_858 ,
       \genblk1[12].inst_SUB_UNS_OP_n_859 ,
       \genblk1[12].inst_SUB_UNS_OP_n_862 ,
       \genblk1[12].inst_SUB_UNS_OP_n_865 ;
  wire \genblk1[12].inst_SUB_UNS_OP_n_866 ,
       \genblk1[12].inst_SUB_UNS_OP_n_867 ,
       \genblk1[12].inst_SUB_UNS_OP_n_869 ,
       \genblk1[12].inst_SUB_UNS_OP_n_871 ,
       \genblk1[12].inst_SUB_UNS_OP_n_873 ,
       \genblk1[12].inst_SUB_UNS_OP_n_874 ,
       \genblk1[12].inst_SUB_UNS_OP_n_876 , \genblk1[12].inst_n_709 ;
  wire \genblk1[12].inst_n_710 , \genblk1[12].inst_n_711 ,
       \genblk1[12].inst_n_712 , \genblk1[12].inst_n_713 ,
       \genblk1[12].inst_n_714 , \genblk1[12].inst_n_715 ,
       \genblk1[12].inst_n_716 , \genblk1[12].inst_n_717 ;
  wire \genblk1[12].inst_n_718 , \genblk1[12].inst_n_719 ,
       \genblk1[13].inst_SUB_UNS_OP_n_869 ,
       \genblk1[13].inst_SUB_UNS_OP_n_872 ,
       \genblk1[13].inst_SUB_UNS_OP_n_874 ,
       \genblk1[13].inst_SUB_UNS_OP_n_876 ,
       \genblk1[13].inst_SUB_UNS_OP_n_878 ,
       \genblk1[13].inst_SUB_UNS_OP_n_880 ;
  wire \genblk1[13].inst_SUB_UNS_OP_n_882 ,
       \genblk1[13].inst_SUB_UNS_OP_n_884 ,
       \genblk1[13].inst_SUB_UNS_OP_n_886 ,
       \genblk1[13].inst_SUB_UNS_OP_n_888 ,
       \genblk1[13].inst_SUB_UNS_OP_n_890 ,
       \genblk1[13].inst_SUB_UNS_OP_n_892 ,
       \genblk1[13].inst_SUB_UNS_OP_n_894 ,
       \genblk1[13].inst_SUB_UNS_OP_n_895 ;
  wire \genblk1[13].inst_SUB_UNS_OP_n_896 ,
       \genblk1[13].inst_SUB_UNS_OP_n_898 ,
       \genblk1[13].inst_SUB_UNS_OP_n_899 ,
       \genblk1[13].inst_SUB_UNS_OP_n_901 ,
       \genblk1[13].inst_SUB_UNS_OP_n_902 ,
       \genblk1[13].inst_SUB_UNS_OP_n_903 ,
       \genblk1[13].inst_SUB_UNS_OP_n_904 ,
       \genblk1[13].inst_SUB_UNS_OP_n_905 ;
  wire \genblk1[13].inst_SUB_UNS_OP_n_906 ,
       \genblk1[13].inst_SUB_UNS_OP_n_907 ,
       \genblk1[13].inst_SUB_UNS_OP_n_911 ,
       \genblk1[13].inst_SUB_UNS_OP_n_916 ,
       \genblk1[13].inst_SUB_UNS_OP_n_919 ,
       \genblk1[13].inst_SUB_UNS_OP_n_920 ,
       \genblk1[13].inst_SUB_UNS_OP_n_921 ,
       \genblk1[13].inst_SUB_UNS_OP_n_923 ;
  wire \genblk1[13].inst_SUB_UNS_OP_n_924 ,
       \genblk1[13].inst_SUB_UNS_OP_n_927 , \genblk1[13].inst_n_710 ,
       \genblk1[13].inst_n_711 , \genblk1[13].inst_n_712 ,
       \genblk1[13].inst_n_713 , \genblk1[13].inst_n_714 ,
       \genblk1[13].inst_n_715 ;
  wire \genblk1[13].inst_n_716 , \genblk1[13].inst_n_717 ,
       \genblk1[13].inst_n_718 , \genblk1[13].inst_n_719 ,
       \genblk1[13].inst_n_720 , \genblk1[13].inst_n_721 ,
       \genblk1[14].inst_SUB_UNS_OP_n_909 ,
       \genblk1[14].inst_SUB_UNS_OP_n_912 ;
  wire \genblk1[14].inst_SUB_UNS_OP_n_914 ,
       \genblk1[14].inst_SUB_UNS_OP_n_916 ,
       \genblk1[14].inst_SUB_UNS_OP_n_918 ,
       \genblk1[14].inst_SUB_UNS_OP_n_920 ,
       \genblk1[14].inst_SUB_UNS_OP_n_922 ,
       \genblk1[14].inst_SUB_UNS_OP_n_924 ,
       \genblk1[14].inst_SUB_UNS_OP_n_926 ,
       \genblk1[14].inst_SUB_UNS_OP_n_928 ;
  wire \genblk1[14].inst_SUB_UNS_OP_n_930 ,
       \genblk1[14].inst_SUB_UNS_OP_n_932 ,
       \genblk1[14].inst_SUB_UNS_OP_n_934 ,
       \genblk1[14].inst_SUB_UNS_OP_n_935 ,
       \genblk1[14].inst_SUB_UNS_OP_n_936 ,
       \genblk1[14].inst_SUB_UNS_OP_n_938 ,
       \genblk1[14].inst_SUB_UNS_OP_n_939 ,
       \genblk1[14].inst_SUB_UNS_OP_n_940 ;
  wire \genblk1[14].inst_SUB_UNS_OP_n_941 ,
       \genblk1[14].inst_SUB_UNS_OP_n_943 ,
       \genblk1[14].inst_SUB_UNS_OP_n_945 ,
       \genblk1[14].inst_SUB_UNS_OP_n_947 ,
       \genblk1[14].inst_SUB_UNS_OP_n_949 ,
       \genblk1[14].inst_SUB_UNS_OP_n_950 ,
       \genblk1[14].inst_SUB_UNS_OP_n_951 ,
       \genblk1[14].inst_SUB_UNS_OP_n_952 ;
  wire \genblk1[14].inst_SUB_UNS_OP_n_953 ,
       \genblk1[14].inst_SUB_UNS_OP_n_955 ,
       \genblk1[14].inst_SUB_UNS_OP_n_956 ,
       \genblk1[14].inst_SUB_UNS_OP_n_959 ,
       \genblk1[14].inst_SUB_UNS_OP_n_960 ,
       \genblk1[14].inst_SUB_UNS_OP_n_961 ,
       \genblk1[14].inst_SUB_UNS_OP_n_964 ,
       \genblk1[14].inst_SUB_UNS_OP_n_966 ;
  wire \genblk1[14].inst_SUB_UNS_OP_n_968 ,
       \genblk1[14].inst_SUB_UNS_OP_n_972 , \genblk1[14].inst_n_711 ,
       \genblk1[14].inst_n_712 , \genblk1[14].inst_n_713 ,
       \genblk1[14].inst_n_714 , \genblk1[14].inst_n_715 ,
       \genblk1[14].inst_n_716 ;
  wire \genblk1[14].inst_n_717 , \genblk1[14].inst_n_718 ,
       \genblk1[14].inst_n_719 , \genblk1[14].inst_n_720 ,
       \genblk1[14].inst_n_721 , \genblk1[14].inst_n_722 ,
       \genblk1[14].inst_n_723 , \genblk1[15].inst_SUB_UNS_OP_n_893 ;
  wire \genblk1[15].inst_SUB_UNS_OP_n_898 ,
       \genblk1[15].inst_SUB_UNS_OP_n_909 ,
       \genblk1[15].inst_SUB_UNS_OP_n_911 ,
       \genblk1[15].inst_SUB_UNS_OP_n_941 ,
       \genblk1[15].inst_SUB_UNS_OP_n_943 ,
       \genblk1[15].inst_SUB_UNS_OP_n_948 ,
       \genblk1[15].inst_SUB_UNS_OP_n_949 ,
       \genblk1[15].inst_SUB_UNS_OP_n_954 ;
  wire \genblk1[15].inst_SUB_UNS_OP_n_957 ,
       \genblk1[15].inst_SUB_UNS_OP_n_959 ,
       \genblk1[15].inst_SUB_UNS_OP_n_961 ,
       \genblk1[15].inst_SUB_UNS_OP_n_963 ,
       \genblk1[15].inst_SUB_UNS_OP_n_965 ,
       \genblk1[15].inst_SUB_UNS_OP_n_967 ,
       \genblk1[15].inst_SUB_UNS_OP_n_969 ,
       \genblk1[15].inst_SUB_UNS_OP_n_971 ;
  wire \genblk1[15].inst_SUB_UNS_OP_n_973 ,
       \genblk1[15].inst_SUB_UNS_OP_n_975 ,
       \genblk1[15].inst_SUB_UNS_OP_n_977 ,
       \genblk1[15].inst_SUB_UNS_OP_n_979 ,
       \genblk1[15].inst_SUB_UNS_OP_n_981 ,
       \genblk1[15].inst_SUB_UNS_OP_n_983 ,
       \genblk1[15].inst_SUB_UNS_OP_n_984 ,
       \genblk1[15].inst_SUB_UNS_OP_n_985 ;
  wire \genblk1[15].inst_SUB_UNS_OP_n_987 ,
       \genblk1[15].inst_SUB_UNS_OP_n_988 ,
       \genblk1[15].inst_SUB_UNS_OP_n_990 ,
       \genblk1[15].inst_SUB_UNS_OP_n_991 ,
       \genblk1[15].inst_SUB_UNS_OP_n_992 ,
       \genblk1[15].inst_SUB_UNS_OP_n_993 ,
       \genblk1[15].inst_SUB_UNS_OP_n_994 ,
       \genblk1[15].inst_SUB_UNS_OP_n_998 ;
  wire \genblk1[15].inst_SUB_UNS_OP_n_999 ,
       \genblk1[15].inst_SUB_UNS_OP_n_1004 ,
       \genblk1[15].inst_SUB_UNS_OP_n_1007 ,
       \genblk1[15].inst_SUB_UNS_OP_n_1008 ,
       \genblk1[15].inst_SUB_UNS_OP_n_1011 ,
       \genblk1[15].inst_SUB_UNS_OP_n_1012 ,
       \genblk1[15].inst_SUB_UNS_OP_n_1016 ,
       \genblk1[15].inst_SUB_UNS_OP_n_1017 ;
  wire \genblk1[15].inst_SUB_UNS_OP_n_1018 ,
       \genblk1[15].inst_SUB_UNS_OP_n_1019 ,
       \genblk1[15].inst_SUB_UNS_OP_n_1026 ,
       \genblk1[15].inst_SUB_UNS_OP_n_1028 ,
       \genblk1[15].inst_SUB_UNS_OP_n_1029 ,
       \genblk1[15].inst_SUB_UNS_OP_n_1030 ,
       \genblk1[15].inst_SUB_UNS_OP_n_1031 ,
       \genblk1[15].inst_SUB_UNS_OP_n_1032 ;
  wire \genblk1[15].inst_SUB_UNS_OP_n_1033 ,
       \genblk1[15].inst_SUB_UNS_OP_n_1034 , \genblk1[15].inst_n_712 ,
       \genblk1[15].inst_n_713 , \genblk1[15].inst_n_714 ,
       \genblk1[15].inst_n_715 , \genblk1[15].inst_n_716 ,
       \genblk1[15].inst_n_717 ;
  wire \genblk1[15].inst_n_718 , \genblk1[15].inst_n_719 ,
       \genblk1[15].inst_n_720 , \genblk1[15].inst_n_721 ,
       \genblk1[15].inst_n_722 , \genblk1[15].inst_n_723 ,
       \genblk1[15].inst_n_724 , \genblk1[15].inst_n_725 ;
  wire \genblk1[15].inst_n_1114 , n_0, n_1, n_2, n_3, n_4, n_5, n_6;
  wire n_7, n_8, n_9, n_10, n_11, n_12, n_13, n_14;
  wire n_15, n_16, n_17, n_18, n_19, n_20, n_21, n_22;
  wire n_23, n_24, n_25, n_26, n_27, n_28, n_29, n_30;
  wire n_31, n_32, n_33, n_34, n_35, n_36, n_37, n_38;
  wire n_39, n_40, n_41, n_42, n_43, n_44, n_45, n_46;
  wire n_47, n_48, n_49, n_50, n_51, n_52, n_53, n_54;
  wire n_55, n_56, n_57, n_58, n_59, n_60, n_61, n_62;
  wire n_63, n_64, n_65, n_66, n_67, n_68, n_69, n_70;
  wire n_71, n_72, n_73, n_74, n_75, n_76, n_77, n_78;
  wire n_79, n_80, n_81, n_82, n_83, n_84, n_85, n_86;
  wire n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94;
  wire n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102;
  wire n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110;
  wire n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118;
  wire n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158;
  wire n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166;
  wire n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174;
  wire n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182;
  wire n_183, n_184, n_185, n_186, n_187, n_188, n_189, n_190;
  wire n_191, n_192, n_193, n_194, n_195, n_196, n_197, n_198;
  wire n_199, n_200, n_201, n_202, n_203, n_204, n_205, n_206;
  wire n_207, n_208, n_209, n_210, n_211, n_212, n_213, n_214;
  wire n_215, n_216, n_217, n_218, n_219, n_220, n_221, n_222;
  wire n_223, n_224, n_225, n_226, n_227, n_228, n_229, n_230;
  wire n_231, n_232, n_233, n_234, n_235, n_236, n_237, n_238;
  wire n_239, n_240, n_241, n_242, n_243, n_244, n_245, n_246;
  wire n_247, n_248, n_249, n_250, n_251, n_252, n_253, n_254;
  wire n_255, n_256, n_257, n_258, n_259, n_260, n_261, n_262;
  wire n_263, n_264, n_265, n_266, n_267, n_268, n_269, n_270;
  wire n_271, n_272, n_273, n_274, n_275, n_276, n_277, n_278;
  wire n_279, n_280, n_281, n_282, n_283, n_284, n_285, n_286;
  wire n_287, n_288, n_289, n_290, n_291, n_292, n_293, n_294;
  wire n_295, n_296, n_297, n_298, n_299, n_300, n_301, n_302;
  wire n_303, n_304, n_305, n_306, n_307, n_308, n_309, n_310;
  wire n_311, n_312, n_313, n_314, n_315, n_316, n_317, n_318;
  wire n_319, n_320, n_321, n_322, n_323, n_324, n_325, n_326;
  wire n_327, n_328, n_329, n_330, n_331, n_332, n_333, n_334;
  wire n_335, n_336, n_337, n_338, n_339, n_340, n_341, n_342;
  wire n_343, n_344, n_345, n_346, n_347, n_348, n_349, n_350;
  wire n_351, n_352, n_353, n_354, n_355, n_356, n_357, n_358;
  wire n_359, n_360, n_361, n_362, n_363, n_364, n_365, n_366;
  wire n_367, n_368, n_369, n_370, n_371, n_372, n_373, n_374;
  wire n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382;
  wire n_383, n_384, n_385, n_386, n_387, n_388, n_389, n_390;
  wire n_391, n_392, n_393, n_394, n_395, n_396, n_397, n_398;
  wire n_399, n_400, n_401, n_402, n_403, n_404, n_405, n_406;
  wire n_407, n_408, n_409, n_410, n_411, n_412, n_413, n_414;
  wire n_415, n_416, n_417, n_418, n_419, n_420, n_421, n_422;
  wire n_423, n_424, n_425, n_426, n_427, n_428, n_429, n_430;
  wire n_431, n_432, n_433, n_434, n_435, n_436, n_437, n_438;
  wire n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446;
  wire n_447, n_448, n_449, n_450, n_451, n_452, n_453, n_454;
  wire n_455, n_456, n_457, n_458, n_459, n_460, n_461, n_462;
  wire n_463, n_464, n_465, n_466, n_467, n_468, n_469, n_470;
  wire n_471, n_472, n_473, n_474, n_475, n_476, n_477, n_478;
  wire n_479, n_480, n_481, n_482, n_483, n_484, n_485, n_486;
  wire n_487, n_488, n_489, n_490, n_491, n_492, n_493, n_494;
  wire n_495, n_496, n_497, n_498, n_499, n_500, n_501, n_502;
  wire n_503, n_504, n_505, n_506, n_507, n_508, n_509, n_510;
  wire n_511, n_512, n_513, n_514, n_515, n_516, n_517, n_518;
  wire n_519, n_520, n_521, n_522, n_523, n_524, n_525, n_526;
  wire n_527, n_528, n_529, n_530, n_531, n_532, n_533, n_534;
  wire n_535, n_536, n_537, n_538, n_539, n_540, n_541, n_542;
  wire n_543, n_544, n_545, n_546, n_547, n_548, n_549, n_550;
  wire n_551, n_552, n_553, n_554, n_555, n_556, n_557, n_558;
  wire n_559, n_560, n_561, n_562, n_563, n_564, n_565, n_566;
  wire n_567, n_568, n_569, n_570, n_571, n_572, n_573, n_574;
  wire n_575, n_576, n_577, n_578, n_579, n_580, n_581, n_582;
  wire n_583, n_584, n_585, n_586, n_587, n_588, n_589, n_590;
  wire n_591, n_592, n_593, n_594, n_595, n_596, n_597, n_598;
  wire n_599, n_600, n_601, n_602, n_603, n_604, n_605, n_606;
  wire n_607, n_608, n_609, n_610, n_611, n_612, n_613, n_614;
  wire n_615, n_616, n_617, n_618, n_619, n_620, n_621, n_622;
  wire n_623, n_624, n_625, n_626, n_627, n_628, n_629, n_630;
  wire n_631, n_632, n_633, n_634, n_635, n_636, n_637, n_638;
  wire n_639, n_640, n_641, n_642, n_643, n_644, n_645, n_646;
  wire n_647, n_648, n_649, n_650, n_651, n_652, n_653, n_654;
  wire n_655, n_656, n_657, n_658, n_659, n_660, n_661, n_662;
  wire n_663, n_664, n_665, n_666, n_667, n_668, n_669, n_670;
  wire n_671, n_672, n_673, n_674, n_675, n_676, n_677, n_678;
  wire n_679, n_680, n_681, n_682, n_683, n_684, n_685, n_686;
  wire n_687, n_688, n_689, n_690, n_691, n_692, n_693, n_694;
  wire n_695, n_696, n_697, n_698, n_699, n_700, n_701, n_702;
  wire n_703, n_704, n_705, n_706, n_707, n_708, n_709, n_710;
  wire n_711, n_712, n_713, n_714, n_715, n_716, n_717, n_718;
  wire n_719, n_720, n_721, n_722, n_723, n_724, n_725, n_726;
  wire n_727, n_728, n_729, n_730, n_731, n_732, n_733, n_734;
  wire n_735, n_736, n_737, n_738, n_739, n_740, n_741, n_742;
  wire n_743, n_744, n_745, n_746, n_747, n_748, n_749, n_750;
  wire n_751, n_752, n_753, n_754, n_755, n_756, n_757, n_758;
  wire n_759, n_760, n_761, n_762, n_763, n_764, n_765, n_766;
  wire n_767, n_768, n_769, n_770, n_771, n_772, n_773, n_774;
  wire n_775, n_776, n_777, n_778, n_779, n_780, n_781, n_782;
  wire n_783, n_784, n_785, n_786, n_787, n_788, n_789, n_790;
  wire n_791, n_792, n_793, n_794, n_795, n_796, n_797, n_798;
  wire n_799, n_800, n_801, n_802, n_803, n_804, n_805, n_806;
  wire n_807, n_808, n_809, n_810, n_811, n_812, n_813, n_814;
  wire n_815, n_816, n_817, n_818, n_819, n_820, n_821, n_822;
  wire n_823, n_824, n_825, n_826, n_827, n_828, n_829, n_830;
  wire n_831, n_832, n_833, n_834, n_835, n_836, n_837, n_838;
  wire n_839, n_840, n_841, n_842, n_843, n_844, n_845, n_846;
  wire n_847, n_848, n_849, n_850, n_851, n_852, n_853, n_854;
  wire n_855, n_856, n_857, n_858, n_859, n_860, n_861, n_862;
  wire n_863, n_864, n_865, n_866, n_867, n_868, n_869, n_870;
  wire n_871, n_872, n_873, n_874, n_875, n_876, n_877, n_878;
  wire n_879, n_880, n_881, n_882, n_883, n_884, n_885, n_886;
  wire n_887, n_888, n_889, n_890, n_891, n_892, n_893, n_894;
  wire n_895, n_896, n_897, n_898, n_899, n_900, n_901, n_902;
  wire n_903, n_904, n_905, n_906, n_907, n_908, n_909, n_910;
  wire n_911, n_912, n_913, n_914, n_915, n_916, n_917, n_918;
  wire n_919, n_920, n_921, n_922, n_923, n_924, n_925, n_926;
  wire n_927, n_928, n_929, n_930, n_931, n_932, n_933, n_934;
  wire n_935, n_936, n_937, n_938, n_939, n_940, n_941, n_942;
  wire n_943, n_944, n_945, n_946, n_947, n_948, n_949, n_950;
  wire n_951, n_952, n_953, n_954, n_955, n_956, n_957, n_958;
  wire n_959, n_960, n_961, n_962, n_963, n_964, n_965, n_966;
  wire n_967, n_968, n_969, n_970, n_971, n_972, n_973, n_974;
  wire n_975, n_976, n_977, n_978, n_979, n_980, n_981, n_982;
  wire n_983, n_984, n_985, n_986, n_987, n_988, n_989, n_990;
  wire n_991, n_992, n_993, n_994, n_995;
  NOR2X1 g3518(.A (\genblk1[15].inst_n_1114 ), .B (n_994), .Y (n_995));
  AND2X1 g3519(.A (result[2]), .B (result[15]), .Y
       (\genblk1[14].inst_n_711 ));
  AND2X1 g3520(.A (result[2]), .B (result[14]), .Y
       (\genblk1[14].inst_n_712 ));
  AND2X1 g3521(.A (result[2]), .B (result[13]), .Y
       (\genblk1[14].inst_n_713 ));
  AND2X1 g3522(.A (result[2]), .B (result[12]), .Y
       (\genblk1[14].inst_n_714 ));
  AND2X1 g3523(.A (result[2]), .B (result[10]), .Y
       (\genblk1[14].inst_n_716 ));
  AND2X1 g3524(.A (result[2]), .B (result[3]), .Y
       (\genblk1[14].inst_n_723 ));
  AND2X1 g3525(.A (result[2]), .B (result[8]), .Y
       (\genblk1[14].inst_n_718 ));
  AND2X1 g3526(.A (result[2]), .B (result[7]), .Y
       (\genblk1[14].inst_n_719 ));
  AND2X1 g3527(.A (result[2]), .B (result[6]), .Y
       (\genblk1[14].inst_n_720 ));
  AND2X1 g3528(.A (result[2]), .B (result[5]), .Y
       (\genblk1[14].inst_n_721 ));
  AND2X1 g3529(.A (result[2]), .B (result[4]), .Y
       (\genblk1[14].inst_n_722 ));
  AND2X1 g3530(.A (result[2]), .B (result[9]), .Y
       (\genblk1[14].inst_n_717 ));
  INVX1 g3531(.A (result[2]), .Y (n_994));
  OR2X1 g3532(.A (n_914), .B (n_913), .Y (result[2]));
  NAND3X1 g3533(.A (n_992), .B (n_920), .C (n_927), .Y (n_993));
  NOR3X1 g3534(.A (1'b0), .B (1'b0), .C (n_991), .Y (n_992));
  OR2X1 g3535(.A (1'b0), .B (n_907), .Y (n_991));
  NAND2X1 g3536(.A (n_905), .B (n_903), .Y (n_990));
  NOR2X1 g3537(.A (\eps[13] [19]), .B (n_911), .Y (n_989));
  AOI21X1 g3538(.A (n_919), .B (n_967), .C (n_909), .Y (n_988));
  AOI21X1 g3539(.A (n_936), .B (\eps[13] [15]), .C (n_912), .Y (n_987));
  AOI22X1 g3540(.A (n_985), .B (n_923), .C (result[12]), .D (n_940), .Y
       (n_986));
  OAI21X1 g3541(.A (\genblk1[15].inst_n_1114 ), .B (\eps[13] [14]), .C
       (n_904), .Y (n_985));
  AOI22X1 g3542(.A (n_925), .B (n_921), .C (result[10]), .D (n_937), .Y
       (n_984));
  AOI22X1 g3543(.A (n_982), .B (n_956), .C (n_935), .D (\eps[13] [13]),
       .Y (n_983));
  OR2X1 g3544(.A (n_978), .B (n_908), .Y (n_982));
  NAND3X1 g3545(.A (n_968), .B (n_972), .C (n_928), .Y (n_981));
  NAND3X1 g3546(.A (n_955), .B (n_922), .C (n_965), .Y (n_980));
  AOI21X1 g3547(.A (result[5]), .B (n_939), .C (n_906), .Y (n_979));
  OAI21X1 g3548(.A (result[8]), .B (n_938), .C (n_977), .Y (n_978));
  OR2X1 g3549(.A (n_918), .B (result[5]), .Y (n_977));
  AOI21X1 g3550(.A (n_931), .B (\eps[13] [7]), .C (n_910), .Y (n_976));
  NAND3X1 g3551(.A (n_969), .B (n_945), .C (n_926), .Y (n_975));
  AOI22X1 g3552(.A (n_966), .B (\eps[13] [16]), .C (n_930), .D
       (\eps[13] [18]), .Y (n_974));
  NAND2X1 g3553(.A (\eps[13] [8]), .B (n_965), .Y (n_973));
  OR2X1 g3554(.A (n_917), .B (result[6]), .Y (n_972));
  AOI22X1 g3555(.A (n_924), .B (n_941), .C (result[3]), .D (n_944), .Y
       (n_971));
  NAND2X1 g3556(.A (\eps[13] [9]), .B (n_961), .Y (n_970));
  OR2X1 g3557(.A (n_915), .B (result[14]), .Y (n_969));
  OR2X1 g3558(.A (n_916), .B (result[7]), .Y (n_968));
  INVX1 g3559(.A (n_966), .Y (n_967));
  NAND3X1 g3560(.A (\eps[13] [16]), .B (n_957), .C (n_951), .Y (n_964));
  NOR3X1 g3561(.A (result[13]), .B (n_958), .C (n_952), .Y (n_966));
  AND2X1 g3562(.A (n_961), .B (n_954), .Y (n_965));
  NAND2X1 g3563(.A (\eps[13] [10]), .B (n_929), .Y (n_963));
  NAND2X1 g3564(.A (\eps[13] [17]), .B (n_951), .Y (n_962));
  AOI21X1 g3565(.A (n_933), .B (\eps[13] [6]), .C (query[5]), .Y
       (n_960));
  AND2X1 g3566(.A (n_929), .B (n_953), .Y (n_961));
  INVX1 g3567(.A (n_957), .Y (n_958));
  OR2X1 g3568(.A (\eps[13] [12]), .B (n_932), .Y (n_956));
  OR2X1 g3569(.A (\eps[13] [7]), .B (n_931), .Y (n_955));
  OR2X1 g3570(.A (\eps[13] [9]), .B (n_934), .Y (n_954));
  OR2X1 g3571(.A (\eps[13] [10]), .B (n_942), .Y (n_953));
  NAND2X1 g3572(.A (result[8]), .B (n_938), .Y (n_959));
  OR2X1 g3573(.A (\eps[13] [17]), .B (n_943), .Y (n_957));
  INVX1 g3574(.A (n_951), .Y (n_952));
  NOR2X1 g3575(.A (1'b0), .B (1'b0), .Y (n_950));
  NOR2X1 g3576(.A (1'b0), .B (1'b0), .Y (n_949));
  NAND2X1 g3577(.A (n_932), .B (\eps[13] [12]), .Y (n_948));
  NAND2X1 g3578(.A (\genblk1[15].inst_n_1114 ), .B (\eps[13] [14]), .Y
       (n_947));
  NOR2X1 g3579(.A (1'b0), .B (1'b0), .Y (n_946));
  OR2X1 g3580(.A (\eps[13] [18]), .B (n_930), .Y (n_951));
  INVX1 g3581(.A (\eps[13] [24]), .Y (n_945));
  INVX1 g3582(.A (\eps[13] [6]), .Y (n_944));
  INVX1 g3583(.A (result[14]), .Y (n_943));
  INVX1 g3584(.A (result[7]), .Y (n_942));
  INVX1 g3585(.A (query[4]), .Y (n_941));
  INVX1 g3586(.A (\eps[13] [15]), .Y (n_940));
  INVX1 g3587(.A (\eps[13] [8]), .Y (n_939));
  INVX1 g3588(.A (\eps[13] [11]), .Y (n_938));
  INVX1 g3589(.A (\eps[13] [13]), .Y (n_937));
  INVX1 g3590(.A (result[12]), .Y (n_936));
  INVX1 g3591(.A (result[10]), .Y (n_935));
  INVX1 g3592(.A (result[6]), .Y (n_934));
  INVX1 g3593(.A (result[3]), .Y (n_933));
  INVX1 g3594(.A (result[9]), .Y (n_932));
  INVX1 g3595(.A (result[4]), .Y (n_931));
  INVX1 g3596(.A (result[15]), .Y (n_930));
  BUFX2 drc_bufs3600(.A (n_980), .Y (n_928));
  BUFX2 drc_bufs3601(.A (n_950), .Y (n_927));
  BUFX2 drc_bufs3602(.A (n_949), .Y (n_926));
  BUFX2 drc_bufs3603(.A (n_983), .Y (n_925));
  BUFX2 drc_bufs3604(.A (n_960), .Y (n_924));
  BUFX2 drc_bufs3605(.A (n_947), .Y (n_923));
  BUFX2 drc_bufs3606(.A (n_979), .Y (n_922));
  BUFX2 drc_bufs3607(.A (n_948), .Y (n_921));
  BUFX2 drc_bufs3608(.A (n_946), .Y (n_920));
  BUFX2 drc_bufs3609(.A (n_964), .Y (n_919));
  BUFX2 drc_bufs3610(.A (n_973), .Y (n_918));
  BUFX2 drc_bufs3611(.A (n_970), .Y (n_917));
  BUFX2 drc_bufs3612(.A (n_963), .Y (n_916));
  BUFX2 drc_bufs3613(.A (n_962), .Y (n_915));
  BUFX2 drc_bufs3614(.A (n_993), .Y (n_914));
  BUFX2 drc_bufs3615(.A (n_975), .Y (n_913));
  BUFX2 drc_bufs3616(.A (n_986), .Y (n_912));
  BUFX2 drc_bufs3617(.A (n_988), .Y (n_911));
  BUFX2 drc_bufs3618(.A (n_971), .Y (n_910));
  BUFX2 drc_bufs3619(.A (n_987), .Y (n_909));
  BUFX2 drc_bufs3620(.A (n_981), .Y (n_908));
  BUFX2 drc_bufs3621(.A (n_990), .Y (n_907));
  BUFX2 drc_bufs3622(.A (n_976), .Y (n_906));
  BUFX2 drc_bufs3623(.A (n_974), .Y (n_905));
  BUFX2 drc_bufs3624(.A (n_984), .Y (n_904));
  BUFX2 drc_bufs3625(.A (n_989), .Y (n_903));
  BUFX2 drc_bufs3626(.A (n_995), .Y (\genblk1[14].inst_n_715 ));
  BUFX2 drc_bufs3627(.A (n_959), .Y (n_929));
  AND2X1 g12158(.A (result[6]), .B (result[13]), .Y
       (\genblk1[10].inst_n_709 ));
  AND2X1 g12159(.A (result[6]), .B (result[14]), .Y
       (\genblk1[10].inst_n_708 ));
  AND2X1 g12160(.A (result[6]), .B (result[15]), .Y
       (\genblk1[10].inst_n_707 ));
  AND2X1 g12161(.A (result[6]), .B (result[12]), .Y
       (\genblk1[10].inst_n_710 ));
  AND2X1 g12162(.A (result[6]), .B (result[9]), .Y
       (\genblk1[10].inst_n_713 ));
  AND2X1 g12163(.A (result[6]), .B (result[10]), .Y
       (\genblk1[10].inst_n_712 ));
  AND2X1 g12164(.A (result[6]), .B (n_587), .Y (\genblk1[10].inst_n_711
       ));
  AND2X1 g12165(.A (result[6]), .B (result[8]), .Y
       (\genblk1[10].inst_n_714 ));
  AND2X1 g12166(.A (result[6]), .B (result[7]), .Y
       (\genblk1[10].inst_n_715 ));
  OR2X1 g12167(.A (n_902), .B (\eps[9] [23]), .Y (result[6]));
  OAI21X1 g12168(.A (result[10]), .B (n_449), .C (n_407), .Y (n_902));
  AOI21X1 g12169(.A (n_497), .B (\eps[9] [22]), .C (n_900), .Y (n_901));
  OAI21X1 g12170(.A (n_442), .B (n_898), .C (n_408), .Y (n_900));
  NAND2X1 g12171(.A (\eps[9] [17]), .B (n_896), .Y (n_899));
  OAI21X1 g12172(.A (n_638), .B (\eps[9] [17]), .C (n_896), .Y (n_898));
  AOI21X1 g12173(.A (n_892), .B (n_893), .C (n_433), .Y (n_897));
  AND2X1 g12174(.A (n_484), .B (n_877), .Y (n_896));
  NOR2X1 g12175(.A (n_413), .B (n_458), .Y (n_895));
  NAND3X1 g12177(.A (n_884), .B (n_887), .C (n_893), .Y (n_894));
  XNOR2X1 g12178(.A (n_891), .B (n_392), .Y (\eps[9] [23]));
  OR2X1 g12179(.A (\eps[9] [22]), .B (n_497), .Y (n_893));
  OAI21X1 g12180(.A (result[14]), .B (n_885), .C (n_404), .Y (n_892));
  AND2X1 g12181(.A (n_417), .B (n_857), .Y (n_891));
  NAND3X1 g12182(.A (n_518), .B (\eps[9] [20]), .C (n_887), .Y (n_890));
  XNOR2X1 g12183(.A (n_888), .B (n_859), .Y (\eps[9] [22]));
  NAND2X1 g12184(.A (n_850), .B (n_888), .Y (n_889));
  OR2X1 g12185(.A (n_886), .B (n_843), .Y (n_888));
  OR2X1 g12186(.A (\eps[9] [21]), .B (n_504), .Y (n_887));
  OAI21X1 g12187(.A (n_482), .B (n_882), .C (n_813), .Y (n_886));
  INVX1 g12188(.A (\eps[9] [21]), .Y (n_885));
  AND2X1 g12189(.A (n_883), .B (n_880), .Y (n_884));
  XOR2X1 g12190(.A (n_882), .B (n_863), .Y (\eps[9] [21]));
  OR2X1 g12191(.A (\eps[9] [20]), .B (n_518), .Y (n_883));
  AND2X1 g12192(.A (n_426), .B (n_854), .Y (n_882));
  AOI22X1 g12193(.A (\eps[9] [18]), .B (\genblk1[15].inst_n_1114 ), .C
       (n_546), .D (\eps[9] [19]), .Y (n_881));
  XNOR2X1 g12194(.A (n_878), .B (n_861), .Y (\eps[9] [20]));
  OR2X1 g12195(.A (\eps[9] [19]), .B (n_546), .Y (n_880));
  NAND2X1 g12196(.A (n_851), .B (n_878), .Y (n_879));
  OAI21X1 g12197(.A (n_439), .B (n_876), .C (n_856), .Y (n_878));
  XOR2X1 g12198(.A (n_876), .B (n_858), .Y (\eps[9] [19]));
  OR2X1 g12199(.A (\eps[9] [18]), .B (\genblk1[15].inst_n_1114 ), .Y
       (n_877));
  AND2X1 g12200(.A (n_425), .B (n_855), .Y (n_876));
  XNOR2X1 g12201(.A (n_873), .B (n_862), .Y (\eps[9] [18]));
  NAND2X1 g12202(.A (n_849), .B (n_873), .Y (n_875));
  AOI22X1 g12203(.A (n_444), .B (n_867), .C (n_692), .D (\eps[9] [16]),
       .Y (n_874));
  OR2X1 g12204(.A (n_872), .B (n_843), .Y (n_873));
  OAI21X1 g12205(.A (n_794), .B (n_868), .C (n_793), .Y (n_872));
  AOI21X1 g12206(.A (result[9]), .B (n_869), .C (n_432), .Y (n_871));
  MUX2X1 g12207(.A (n_483), .B (n_868), .S (n_860), .Y (\eps[9] [17]));
  AOI22X1 g12208(.A (\eps[9] [15]), .B (n_766), .C (n_450), .D (n_866),
       .Y (n_870));
  INVX1 g12209(.A (\eps[9] [16]), .Y (n_869));
  INVX1 g12211(.A (n_483), .Y (n_868));
  FAX1 g12212(.A (n_777), .B (n_844), .C (n_847), .YC (n_483), .YS
       (\eps[9] [16]));
  OR2X1 g12213(.A (\eps[9] [15]), .B (n_766), .Y (n_867));
  OAI21X1 g12214(.A (n_487), .B (n_864), .C (n_847), .Y (\eps[9] [15]));
  OAI21X1 g12215(.A (n_466), .B (result[7]), .C (n_865), .Y (n_866));
  INVX1 g12216(.A (n_865), .Y (\eps[9] [14]));
  HAX1 g12217(.A (n_493), .B (result[7]), .YC (n_864), .YS (n_865));
  OR2X1 g12218(.A (n_852), .B (n_812), .Y (n_863));
  OAI21X1 g12219(.A (n_798), .B (n_843), .C (n_855), .Y (n_862));
  OAI21X1 g12220(.A (n_807), .B (n_843), .C (n_854), .Y (n_861));
  AND2X1 g12221(.A (n_853), .B (n_793), .Y (n_860));
  OAI21X1 g12222(.A (n_820), .B (n_843), .C (n_857), .Y (n_859));
  OAI21X1 g12223(.A (n_802), .B (n_843), .C (n_856), .Y (n_858));
  OAI21X1 g12225(.A (n_504), .B (n_843), .C (n_817), .Y (n_857));
  OAI21X1 g12226(.A (\genblk1[15].inst_n_1114 ), .B (n_843), .C
       (n_800), .Y (n_856));
  OAI21X1 g12227(.A (n_638), .B (n_843), .C (n_796), .Y (n_855));
  MUX2X1 g12228(.A (n_794), .B (n_792), .S (result[7]), .Y (n_853));
  MUX2X1 g12229(.A (n_809), .B (n_811), .S (n_843), .Y (n_852));
  OAI21X1 g12230(.A (n_546), .B (n_843), .C (n_805), .Y (n_854));
  OR2X1 g12231(.A (n_843), .B (n_807), .Y (n_851));
  OR2X1 g12232(.A (n_843), .B (n_820), .Y (n_850));
  OR2X1 g12233(.A (n_843), .B (n_798), .Y (n_849));
  NOR2X1 g12234(.A (n_802), .B (n_843), .Y (n_848));
  NAND2X1 g12235(.A (n_466), .B (result[7]), .Y (n_846));
  OR2X1 g12236(.A (n_843), .B (n_497), .Y (n_845));
  OR2X1 g12237(.A (n_843), .B (n_766), .Y (n_844));
  OR2X1 g12238(.A (n_843), .B (n_501), .Y (n_847));
  INVX1 g12239(.A (result[7]), .Y (n_843));
  OR2X1 g12240(.A (n_842), .B (n_831), .Y (result[7]));
  OAI21X1 g12241(.A (n_784), .B (n_825), .C (n_841), .Y (n_842));
  AND2X1 g12242(.A (n_429), .B (n_422), .Y (n_841));
  AOI22X1 g12243(.A (n_825), .B (n_784), .C (n_501), .D (n_838), .Y
       (n_840));
  AOI21X1 g12244(.A (query[16]), .B (n_837), .C (n_835), .Y (n_839));
  OAI21X1 g12245(.A (n_788), .B (n_834), .C (n_836), .Y (n_838));
  INVX1 g12246(.A (n_836), .Y (n_837));
  OR2X1 g12247(.A (n_834), .B (result[8]), .Y (n_836));
  OAI21X1 g12248(.A (n_793), .B (n_833), .C (n_832), .Y (n_835));
  OR2X1 g12249(.A (n_833), .B (n_794), .Y (n_834));
  OR2X1 g12250(.A (n_830), .B (n_799), .Y (n_833));
  OR2X1 g12251(.A (n_830), .B (n_434), .Y (n_832));
  OAI21X1 g12252(.A (n_506), .B (n_447), .C (n_829), .Y (n_831));
  OR2X1 g12253(.A (n_437), .B (n_482), .Y (n_830));
  OAI21X1 g12254(.A (n_812), .B (n_818), .C (n_826), .Y (n_829));
  NAND3X1 g12255(.A (n_802), .B (n_807), .C (n_826), .Y (n_828));
  AOI22X1 g12256(.A (n_824), .B (n_817), .C (n_497), .D (n_821), .Y
       (n_827));
  AND2X1 g12257(.A (n_823), .B (n_820), .Y (n_826));
  OR2X1 g12258(.A (n_822), .B (n_766), .Y (n_825));
  OR2X1 g12259(.A (n_821), .B (n_505), .Y (n_824));
  OR2X1 g12260(.A (n_821), .B (n_497), .Y (n_823));
  OAI21X1 g12261(.A (n_481), .B (n_819), .C (n_745), .Y (n_822));
  XOR2X1 g12263(.A (n_819), .B (n_787), .Y (n_821));
  OR2X1 g12264(.A (n_817), .B (n_504), .Y (n_820));
  AND2X1 g12265(.A (n_431), .B (n_780), .Y (n_819));
  INVX1 g12266(.A (n_395), .Y (n_818));
  NAND3X1 g12267(.A (n_546), .B (n_805), .C (n_811), .Y (n_816));
  XNOR2X1 g12268(.A (n_814), .B (n_785), .Y (n_817));
  NAND2X1 g12269(.A (n_772), .B (n_814), .Y (n_815));
  OR2X1 g12270(.A (n_810), .B (n_766), .Y (n_814));
  INVX1 g12271(.A (n_812), .Y (n_813));
  INVX1 g12273(.A (n_811), .Y (n_482));
  AND2X1 g12274(.A (n_808), .B (n_518), .Y (n_812));
  OR2X1 g12275(.A (n_808), .B (n_518), .Y (n_811));
  OAI21X1 g12276(.A (n_730), .B (n_806), .C (n_731), .Y (n_810));
  INVX1 g12277(.A (n_808), .Y (n_809));
  XOR2X1 g12278(.A (n_806), .B (n_786), .Y (n_808));
  OR2X1 g12279(.A (n_805), .B (n_546), .Y (n_807));
  AND2X1 g12280(.A (n_421), .B (n_779), .Y (n_806));
  AOI22X1 g12281(.A (n_796), .B (n_638), .C (\genblk1[15].inst_n_1114
       ), .D (n_800), .Y (n_804));
  XNOR2X1 g12282(.A (n_801), .B (n_781), .Y (n_805));
  NAND2X1 g12283(.A (n_771), .B (n_801), .Y (n_803));
  OR2X1 g12284(.A (n_800), .B (\genblk1[15].inst_n_1114 ), .Y (n_802));
  OAI21X1 g12285(.A (n_769), .B (n_797), .C (n_778), .Y (n_801));
  XNOR2X1 g12286(.A (n_797), .B (n_782), .Y (n_800));
  INVX1 g12287(.A (n_798), .Y (n_799));
  OR2X1 g12288(.A (n_796), .B (n_638), .Y (n_798));
  AND2X1 g12289(.A (n_419), .B (n_776), .Y (n_797));
  XNOR2X1 g12290(.A (n_790), .B (n_783), .Y (n_796));
  NAND2X1 g12291(.A (n_767), .B (n_790), .Y (n_795));
  AND2X1 g12292(.A (n_791), .B (result[9]), .Y (n_794));
  OR2X1 g12293(.A (n_791), .B (result[9]), .Y (n_793));
  INVX1 g12294(.A (n_791), .Y (n_792));
  AND2X1 g12295(.A (n_790), .B (n_430), .Y (n_791));
  OR2X1 g12296(.A (n_768), .B (query[17]), .Y (n_790));
  NAND2X1 g12297(.A (query[17]), .B (n_768), .Y (n_789));
  INVX1 g12298(.A (n_777), .Y (n_788));
  OR2X1 g12299(.A (n_775), .B (n_744), .Y (n_787));
  OR2X1 g12300(.A (n_774), .B (n_732), .Y (n_786));
  OAI21X1 g12301(.A (n_738), .B (n_766), .C (n_780), .Y (n_785));
  OAI21X1 g12302(.A (n_479), .B (n_766), .C (n_776), .Y (n_783));
  AND2X1 g12303(.A (n_778), .B (n_770), .Y (n_782));
  OAI21X1 g12304(.A (n_726), .B (n_766), .C (n_779), .Y (n_781));
  OAI21X1 g12305(.A (n_754), .B (n_766), .C (n_773), .Y (n_784));
  OAI21X1 g12306(.A (n_518), .B (n_766), .C (n_736), .Y (n_780));
  OAI21X1 g12307(.A (\genblk1[15].inst_n_1114 ), .B (n_766), .C
       (n_723), .Y (n_779));
  OAI21X1 g12308(.A (n_638), .B (n_766), .C (n_711), .Y (n_778));
  OAI21X1 g12309(.A (n_485), .B (result[8]), .C (n_768), .Y (n_777));
  MUX2X1 g12310(.A (n_740), .B (n_743), .S (n_766), .Y (n_775));
  MUX2X1 g12311(.A (n_728), .B (n_480), .S (n_766), .Y (n_774));
  OAI21X1 g12312(.A (n_497), .B (n_766), .C (n_747), .Y (n_773));
  OAI21X1 g12313(.A (n_692), .B (n_766), .C (n_706), .Y (n_776));
  OR2X1 g12314(.A (n_766), .B (n_738), .Y (n_772));
  OR2X1 g12315(.A (n_766), .B (n_726), .Y (n_771));
  INVX1 g12316(.A (n_769), .Y (n_770));
  OR2X1 g12317(.A (n_766), .B (n_479), .Y (n_767));
  AND2X1 g12318(.A (result[8]), .B (n_720), .Y (n_769));
  OR2X1 g12319(.A (n_766), .B (query[16]), .Y (n_768));
  INVX1 g12320(.A (result[8]), .Y (n_766));
  OR2X1 g12321(.A (n_765), .B (n_756), .Y (result[8]));
  INVX1 g12322(.A (n_397), .Y (n_765));
  AOI22X1 g12323(.A (n_763), .B (n_754), .C (n_712), .D (n_748), .Y
       (n_764));
  OR2X1 g12324(.A (n_762), .B (n_744), .Y (n_763));
  OAI21X1 g12325(.A (n_485), .B (n_760), .C (n_761), .Y (n_762));
  NOR3X1 g12326(.A (n_753), .B (n_454), .C (n_758), .Y (n_761));
  OR2X1 g12327(.A (n_759), .B (n_720), .Y (n_760));
  OR2X1 g12328(.A (n_757), .B (n_708), .Y (n_759));
  NOR3X1 g12329(.A (n_453), .B (n_730), .C (n_755), .Y (n_758));
  OR2X1 g12330(.A (n_755), .B (n_730), .Y (n_757));
  OAI21X1 g12331(.A (n_712), .B (n_748), .C (n_409), .Y (n_756));
  OR2X1 g12332(.A (n_749), .B (n_727), .Y (n_755));
  OR2X1 g12333(.A (n_747), .B (n_497), .Y (n_754));
  INVX1 g12334(.A (n_399), .Y (n_753));
  AOI21X1 g12335(.A (n_731), .B (n_438), .C (n_749), .Y (n_752));
  NAND2X1 g12336(.A (n_497), .B (n_747), .Y (n_751));
  NAND3X1 g12337(.A (n_518), .B (n_736), .C (n_743), .Y (n_750));
  OR2X1 g12338(.A (n_481), .B (n_739), .Y (n_749));
  AND2X1 g12339(.A (n_414), .B (n_709), .Y (n_748));
  XNOR2X1 g12340(.A (n_742), .B (n_714), .Y (n_747));
  NAND2X1 g12341(.A (n_693), .B (n_742), .Y (n_746));
  INVX1 g12342(.A (n_744), .Y (n_745));
  INVX1 g12344(.A (n_743), .Y (n_481));
  AND2X1 g12345(.A (n_741), .B (n_504), .Y (n_744));
  OR2X1 g12346(.A (n_741), .B (n_504), .Y (n_743));
  OAI21X1 g12347(.A (n_700), .B (n_737), .C (n_705), .Y (n_742));
  INVX1 g12348(.A (n_740), .Y (n_741));
  XNOR2X1 g12349(.A (n_737), .B (n_716), .Y (n_740));
  INVX1 g12350(.A (n_738), .Y (n_739));
  OR2X1 g12351(.A (n_736), .B (n_518), .Y (n_738));
  AND2X1 g12352(.A (n_428), .B (n_703), .Y (n_737));
  NAND3X1 g12353(.A (\genblk1[15].inst_n_1114 ), .B (n_723), .C
       (n_480), .Y (n_735));
  XNOR2X1 g12354(.A (n_733), .B (n_715), .Y (n_736));
  NAND2X1 g12355(.A (n_697), .B (n_733), .Y (n_734));
  OR2X1 g12356(.A (n_729), .B (n_692), .Y (n_733));
  INVX1 g12357(.A (n_731), .Y (n_732));
  INVX1 g12359(.A (n_730), .Y (n_480));
  OR2X1 g12360(.A (n_728), .B (result[12]), .Y (n_731));
  AND2X1 g12361(.A (n_728), .B (result[12]), .Y (n_730));
  OAI21X1 g12362(.A (n_474), .B (n_724), .C (n_659), .Y (n_729));
  XNOR2X1 g12363(.A (n_724), .B (n_710), .Y (n_728));
  INVX1 g12364(.A (n_726), .Y (n_727));
  OR2X1 g12365(.A (n_723), .B (\genblk1[15].inst_n_1114 ), .Y (n_726));
  AOI22X1 g12366(.A (n_711), .B (n_638), .C (n_717), .D (n_721), .Y
       (n_725));
  AND2X1 g12367(.A (n_423), .B (n_461), .Y (n_724));
  XNOR2X1 g12368(.A (n_718), .B (n_707), .Y (n_723));
  NAND2X1 g12369(.A (n_695), .B (n_707), .Y (n_722));
  INVX1 g12370(.A (n_720), .Y (n_721));
  AND2X1 g12371(.A (n_719), .B (result[10]), .Y (n_720));
  INVX1 g12372(.A (n_711), .Y (n_719));
  OAI21X1 g12373(.A (n_649), .B (n_692), .C (n_461), .Y (n_718));
  OAI21X1 g12374(.A (n_492), .B (n_708), .C (n_455), .Y (n_717));
  OR2X1 g12375(.A (n_704), .B (n_700), .Y (n_716));
  OAI21X1 g12376(.A (n_663), .B (n_692), .C (n_703), .Y (n_715));
  OAI21X1 g12377(.A (n_679), .B (n_692), .C (n_709), .Y (n_714));
  NAND2X1 g12378(.A (n_649), .B (n_412), .Y (n_713));
  OR2X1 g12379(.A (n_701), .B (n_660), .Y (n_710));
  XNOR2X1 g12380(.A (n_694), .B (n_680), .Y (n_712));
  OAI21X1 g12381(.A (n_495), .B (n_477), .C (n_707), .Y (n_711));
  INVX1 g12383(.A (n_708), .Y (n_479));
  OR2X1 g12384(.A (n_477), .B (n_478), .Y (n_706));
  OAI21X1 g12385(.A (n_504), .B (n_692), .C (n_674), .Y (n_709));
  AND2X1 g12386(.A (n_698), .B (result[9]), .Y (n_708));
  OR2X1 g12387(.A (n_698), .B (query[19]), .Y (n_707));
  INVX1 g12388(.A (n_704), .Y (n_705));
  AOI22X1 g12389(.A (n_642), .B (n_489), .C (result[10]), .D
       (result[9]), .Y (n_702));
  MUX2X1 g12390(.A (n_656), .B (n_658), .S (n_692), .Y (n_701));
  AND2X1 g12391(.A (n_696), .B (n_665), .Y (n_704));
  OAI21X1 g12392(.A (n_546), .B (n_692), .C (n_391), .Y (n_703));
  INVX1 g12395(.A (n_698), .Y (n_477));
  OR2X1 g12396(.A (n_692), .B (n_663), .Y (n_697));
  AND2X1 g12397(.A (result[9]), .B (n_669), .Y (n_700));
  NAND2X1 g12398(.A (query[18]), .B (n_692), .Y (n_699));
  OR2X1 g12399(.A (n_692), .B (query[18]), .Y (n_698));
  OR2X1 g12400(.A (n_692), .B (n_518), .Y (n_696));
  OR2X1 g12401(.A (n_692), .B (n_649), .Y (n_695));
  OR2X1 g12402(.A (n_692), .B (n_497), .Y (n_694));
  OR2X1 g12403(.A (n_692), .B (n_679), .Y (n_693));
  INVX1 g12404(.A (result[9]), .Y (n_692));
  OR2X1 g12405(.A (n_691), .B (n_689), .Y (result[9]));
  OAI21X1 g12406(.A (n_652), .B (n_684), .C (n_411), .Y (n_691));
  AOI22X1 g12407(.A (n_686), .B (n_507), .C (query[18]), .D (n_687), .Y
       (n_690));
  INVX1 g12408(.A (n_398), .Y (n_689));
  AOI22X1 g12409(.A (n_684), .B (n_652), .C (n_682), .D (n_685), .Y
       (n_688));
  AND2X1 g12410(.A (n_685), .B (n_476), .Y (n_687));
  OAI21X1 g12411(.A (n_441), .B (n_680), .C (n_405), .Y (n_686));
  AND2X1 g12412(.A (n_424), .B (n_679), .Y (n_685));
  OR2X1 g12413(.A (n_681), .B (n_638), .Y (n_684));
  NAND2X1 g12414(.A (result[15]), .B (n_680), .Y (n_683));
  OAI21X1 g12415(.A (n_495), .B (n_462), .C (n_403), .Y (n_682));
  OAI21X1 g12416(.A (n_623), .B (n_673), .C (n_624), .Y (n_681));
  MUX2X1 g12417(.A (n_475), .B (n_673), .S (n_460), .Y (n_680));
  NAND2X1 g12418(.A (n_505), .B (n_674), .Y (n_678));
  OR2X1 g12419(.A (n_674), .B (n_504), .Y (n_679));
  NOR2X1 g12421(.A (n_497), .B (n_674), .Y (n_676));
  AOI22X1 g12422(.A (n_672), .B (n_664), .C (n_671), .D (n_668), .Y
       (n_675));
  NAND3X1 g12423(.A (n_649), .B (n_658), .C (n_672), .Y (n_677));
  INVX1 g12425(.A (n_475), .Y (n_673));
  FAX1 g12426(.A (n_613), .B (n_639), .C (n_667), .YC (n_475), .YS
       (n_674));
  AND2X1 g12427(.A (n_668), .B (n_663), .Y (n_672));
  INVX1 g12428(.A (n_396), .Y (n_671));
  AOI22X1 g12429(.A (n_665), .B (n_518), .C (n_546), .D (n_391), .Y
       (n_670));
  INVX1 g12430(.A (n_668), .Y (n_669));
  OR2X1 g12431(.A (n_665), .B (n_518), .Y (n_668));
  INVX1 g12432(.A (n_393), .Y (n_667));
  AOI21X1 g12433(.A (n_644), .B (n_661), .C (n_467), .Y (n_666));
  OAI21X1 g12434(.A (result[10]), .B (n_662), .C (n_659), .Y (n_664));
  XNOR2X1 g12435(.A (n_661), .B (n_653), .Y (n_665));
  OR2X1 g12436(.A (n_391), .B (n_546), .Y (n_663));
  OR2X1 g12437(.A (n_474), .B (n_489), .Y (n_662));
  OAI21X1 g12438(.A (n_440), .B (n_655), .C (n_457), .Y (n_661));
  INVX1 g12440(.A (n_659), .Y (n_660));
  OR2X1 g12441(.A (n_656), .B (n_587), .Y (n_659));
  INVX1 g12443(.A (n_658), .Y (n_474));
  OR2X1 g12444(.A (n_657), .B (\genblk1[15].inst_n_1114 ), .Y (n_658));
  INVX1 g12445(.A (n_656), .Y (n_657));
  HAX1 g12447(.A (n_494), .B (n_641), .YC (n_655), .YS (n_656));
  NAND2X1 g12448(.A (n_624), .B (n_645), .Y (n_654));
  OR2X1 g12449(.A (n_467), .B (n_643), .Y (n_653));
  OAI21X1 g12450(.A (n_592), .B (n_640), .C (n_457), .Y (n_651));
  OAI21X1 g12451(.A (n_630), .B (n_638), .C (n_646), .Y (n_652));
  NAND3X1 g12452(.A (n_599), .B (n_602), .C (n_640), .Y (n_650));
  NOR2X1 g12453(.A (n_592), .B (n_640), .Y (n_648));
  OR2X1 g12454(.A (n_641), .B (n_638), .Y (n_649));
  OAI21X1 g12455(.A (n_497), .B (n_638), .C (n_626), .Y (n_646));
  MUX2X1 g12456(.A (n_623), .B (n_619), .S (result[10]), .Y (n_645));
  AOI21X1 g12457(.A (result[12]), .B (result[10]), .C (n_604), .Y
       (n_647));
  INVX1 g12458(.A (n_643), .Y (n_644));
  INVX1 g12459(.A (n_641), .Y (n_642));
  AND2X1 g12460(.A (result[10]), .B (n_610), .Y (n_643));
  AND2X1 g12461(.A (result[10]), .B (n_489), .Y (n_641));
  OR2X1 g12462(.A (n_638), .B (n_518), .Y (n_639));
  OR2X1 g12463(.A (n_638), .B (\genblk1[15].inst_n_1114 ), .Y (n_640));
  INVX1 g12464(.A (result[10]), .Y (n_638));
  OR2X1 g12465(.A (n_637), .B (n_636), .Y (result[10]));
  OAI21X1 g12466(.A (n_621), .B (n_634), .C (n_402), .Y (n_637));
  OAI21X1 g12467(.A (n_605), .B (n_627), .C (n_401), .Y (n_636));
  AOI22X1 g12468(.A (n_630), .B (n_445), .C (n_605), .D (n_627), .Y
       (n_635));
  OR2X1 g12469(.A (n_632), .B (result[13]), .Y (n_634));
  NAND2X1 g12470(.A (n_624), .B (n_406), .Y (n_633));
  OR2X1 g12471(.A (n_631), .B (n_623), .Y (n_632));
  INVX1 g12472(.A (n_630), .Y (n_631));
  OR2X1 g12473(.A (n_626), .B (n_497), .Y (n_630));
  NAND2X1 g12474(.A (n_497), .B (n_626), .Y (n_629));
  NAND3X1 g12475(.A (n_613), .B (n_616), .C (n_622), .Y (n_628));
  AND2X1 g12476(.A (n_625), .B (n_595), .Y (n_627));
  XOR2X1 g12477(.A (n_620), .B (n_608), .Y (n_626));
  OR2X1 g12478(.A (n_620), .B (n_590), .Y (n_625));
  INVX1 g12479(.A (n_623), .Y (n_622));
  OR2X1 g12480(.A (n_618), .B (result[14]), .Y (n_624));
  AND2X1 g12481(.A (n_618), .B (result[14]), .Y (n_623));
  NOR3X1 g12482(.A (n_611), .B (n_613), .C (n_469), .Y (n_621));
  INVX1 g12483(.A (n_618), .Y (n_619));
  AND2X1 g12484(.A (n_617), .B (n_473), .Y (n_620));
  XNOR2X1 g12485(.A (n_614), .B (n_607), .Y (n_618));
  OR2X1 g12486(.A (n_614), .B (n_593), .Y (n_617));
  OR2X1 g12487(.A (n_469), .B (n_611), .Y (n_616));
  AOI21X1 g12488(.A (n_589), .B (n_603), .C (n_610), .Y (n_615));
  AND2X1 g12489(.A (n_420), .B (n_598), .Y (n_614));
  XNOR2X1 g12490(.A (n_601), .B (n_606), .Y (n_613));
  NAND2X1 g12491(.A (n_588), .B (n_601), .Y (n_612));
  AND2X1 g12492(.A (n_609), .B (n_546), .Y (n_611));
  AND2X1 g12493(.A (n_604), .B (result[12]), .Y (n_610));
  INVX1 g12494(.A (n_604), .Y (n_609));
  OR2X1 g12495(.A (n_596), .B (n_590), .Y (n_608));
  OR2X1 g12496(.A (n_459), .B (n_593), .Y (n_607));
  OAI21X1 g12497(.A (n_562), .B (\genblk1[15].inst_n_1114 ), .C
       (n_598), .Y (n_606));
  OAI21X1 g12498(.A (query[20]), .B (query[21]), .C (n_602), .Y
       (n_603));
  AND2X1 g12499(.A (n_594), .B (n_591), .Y (n_605));
  AND2X1 g12500(.A (n_601), .B (n_416), .Y (n_604));
  NAND2X1 g12501(.A (query[23]), .B (n_472), .Y (n_600));
  OR2X1 g12502(.A (n_592), .B (query[22]), .Y (n_599));
  OR2X1 g12503(.A (n_592), .B (\genblk1[15].inst_n_1114 ), .Y (n_602));
  OR2X1 g12504(.A (n_472), .B (query[23]), .Y (n_601));
  INVX1 g12506(.A (n_595), .Y (n_596));
  OAI21X1 g12507(.A (n_497), .B (\genblk1[15].inst_n_1114 ), .C
       (n_569), .Y (n_594));
  OAI21X1 g12508(.A (n_546), .B (\genblk1[15].inst_n_1114 ), .C
       (n_554), .Y (n_598));
  AOI21X1 g12509(.A (result[13]), .B (n_587), .C (n_559), .Y (n_597));
  OAI21X1 g12510(.A (n_504), .B (\genblk1[15].inst_n_1114 ), .C
       (n_567), .Y (n_595));
  INVX1 g12512(.A (n_592), .Y (n_472));
  OR2X1 g12513(.A (\genblk1[15].inst_n_1114 ), .B (n_575), .Y (n_591));
  AND2X1 g12514(.A (n_587), .B (n_565), .Y (n_593));
  AND2X1 g12515(.A (n_587), .B (n_488), .Y (n_592));
  OR2X1 g12516(.A (n_587), .B (n_488), .Y (n_589));
  AND2X1 g12517(.A (n_587), .B (n_571), .Y (n_590));
  OR2X1 g12518(.A (\genblk1[15].inst_n_1114 ), .B (n_562), .Y (n_588));
  INVX8 g12519(.A (n_587), .Y (\genblk1[15].inst_n_1114 ));
  OAI21X1 g12520(.A (n_563), .B (n_579), .C (n_586), .Y (n_587));
  NOR3X1 g12521(.A (n_581), .B (n_584), .C (n_585), .Y (n_586));
  OAI21X1 g12522(.A (result[13]), .B (n_582), .C (n_580), .Y (n_585));
  OAI21X1 g12523(.A (n_464), .B (n_579), .C (n_583), .Y (n_584));
  OR2X1 g12524(.A (n_436), .B (n_506), .Y (n_583));
  OR2X1 g12525(.A (n_578), .B (n_559), .Y (n_582));
  AND2X1 g12526(.A (n_465), .B (n_560), .Y (n_581));
  OR2X1 g12527(.A (n_465), .B (n_560), .Y (n_580));
  OR2X1 g12528(.A (n_574), .B (n_571), .Y (n_578));
  AOI22X1 g12529(.A (n_569), .B (n_572), .C (n_505), .D (n_567), .Y
       (n_577));
  OR2X1 g12530(.A (n_574), .B (n_573), .Y (n_579));
  NAND3X1 g12531(.A (n_536), .B (result[12]), .C (n_452), .Y (n_576));
  INVX1 g12532(.A (n_574), .Y (n_575));
  OR2X1 g12533(.A (n_571), .B (n_565), .Y (n_573));
  AND2X1 g12534(.A (n_570), .B (result[15]), .Y (n_574));
  OR2X1 g12535(.A (n_567), .B (n_497), .Y (n_572));
  INVX1 g12536(.A (n_569), .Y (n_570));
  AND2X1 g12537(.A (n_566), .B (result[14]), .Y (n_571));
  XNOR2X1 g12538(.A (n_564), .B (n_561), .Y (n_569));
  NAND2X1 g12539(.A (n_534), .B (n_564), .Y (n_568));
  INVX1 g12540(.A (n_566), .Y (n_567));
  XOR2X1 g12541(.A (n_558), .B (n_547), .Y (n_566));
  AND2X1 g12542(.A (n_559), .B (result[13]), .Y (n_565));
  OAI21X1 g12543(.A (query[22]), .B (query[23]), .C (n_562), .Y
       (n_563));
  OAI21X1 g12544(.A (n_548), .B (n_448), .C (n_456), .Y (n_564));
  OR2X1 g12545(.A (n_554), .B (n_546), .Y (n_562));
  OR2X1 g12546(.A (n_552), .B (n_537), .Y (n_561));
  OAI21X1 g12547(.A (n_520), .B (n_549), .C (n_456), .Y (n_558));
  OAI21X1 g12548(.A (n_542), .B (n_546), .C (n_553), .Y (n_560));
  AND2X1 g12549(.A (n_415), .B (n_547), .Y (n_559));
  NAND2X1 g12550(.A (query[25]), .B (n_550), .Y (n_556));
  NOR2X1 g12551(.A (n_520), .B (n_549), .Y (n_555));
  NAND3X1 g12552(.A (n_525), .B (n_523), .C (n_549), .Y (n_557));
  OAI21X1 g12553(.A (n_497), .B (n_546), .C (n_538), .Y (n_553));
  MUX2X1 g12554(.A (n_528), .B (n_534), .S (n_546), .Y (n_552));
  OAI21X1 g12555(.A (query[24]), .B (n_546), .C (n_464), .Y (n_554));
  OR2X1 g12556(.A (n_546), .B (query[24]), .Y (n_550));
  NAND2X1 g12557(.A (query[24]), .B (n_546), .Y (n_551));
  INVX1 g12558(.A (n_547), .Y (n_548));
  OR2X1 g12559(.A (n_546), .B (n_518), .Y (n_549));
  OR2X1 g12560(.A (n_546), .B (n_500), .Y (n_547));
  INVX1 g12561(.A (result[12]), .Y (n_546));
  OR2X1 g12562(.A (n_545), .B (n_543), .Y (result[12]));
  INVX1 g12563(.A (n_394), .Y (n_545));
  AOI22X1 g12564(.A (n_540), .B (n_542), .C (n_468), .D (n_539), .Y
       (n_544));
  OAI21X1 g12565(.A (n_468), .B (n_539), .C (n_410), .Y (n_543));
  OR2X1 g12566(.A (n_538), .B (n_497), .Y (n_542));
  NAND2X1 g12567(.A (n_497), .B (n_538), .Y (n_541));
  OAI21X1 g12568(.A (n_443), .B (n_535), .C (n_536), .Y (n_540));
  AND2X1 g12569(.A (n_418), .B (n_524), .Y (n_539));
  XNOR2X1 g12570(.A (n_527), .B (n_530), .Y (n_538));
  INVX1 g12571(.A (n_536), .Y (n_537));
  OR2X1 g12572(.A (n_528), .B (result[14]), .Y (n_536));
  INVX1 g12573(.A (n_534), .Y (n_535));
  NAND2X1 g12574(.A (n_521), .B (n_527), .Y (n_533));
  OR2X1 g12575(.A (n_532), .B (n_504), .Y (n_534));
  INVX1 g12576(.A (n_528), .Y (n_532));
  AOI22X1 g12577(.A (n_523), .B (n_500), .C (query[26]), .D (n_518), .Y
       (n_531));
  OAI21X1 g12578(.A (n_509), .B (n_519), .C (n_524), .Y (n_530));
  AOI21X1 g12579(.A (n_470), .B (result[13]), .C (n_435), .Y (n_529));
  AND2X1 g12580(.A (n_527), .B (n_427), .Y (n_528));
  AOI21X1 g12581(.A (result[15]), .B (result[13]), .C (n_515), .Y
       (n_526));
  OR2X1 g12582(.A (n_520), .B (query[26]), .Y (n_525));
  OR2X1 g12583(.A (n_471), .B (query[27]), .Y (n_527));
  NAND2X1 g12584(.A (query[27]), .B (n_471), .Y (n_522));
  OAI21X1 g12585(.A (n_508), .B (n_509), .C (n_519), .Y (n_524));
  OR2X1 g12586(.A (n_519), .B (n_509), .Y (n_521));
  OR2X1 g12587(.A (n_520), .B (n_518), .Y (n_523));
  INVX1 g12589(.A (n_520), .Y (n_471));
  AND2X1 g12590(.A (result[13]), .B (n_490), .Y (n_520));
  OR2X1 g12591(.A (n_518), .B (n_504), .Y (n_519));
  INVX1 g12592(.A (result[13]), .Y (n_518));
  OAI21X1 g12593(.A (result[15]), .B (n_515), .C (n_400), .Y
       (result[13]));
  AOI22X1 g12594(.A (n_463), .B (n_446), .C (n_510), .D (n_514), .Y
       (n_517));
  NAND2X1 g12596(.A (result[15]), .B (n_515), .Y (n_516));
  INVX1 g12597(.A (n_513), .Y (n_514));
  HAX1 g12598(.A (n_491), .B (n_509), .YC (n_513), .YS (n_515));
  AOI22X1 g12599(.A (n_511), .B (result[14]), .C (n_490), .D (n_451),
       .Y (n_512));
  INVX1 g12600(.A (n_509), .Y (n_511));
  OAI21X1 g12601(.A (n_502), .B (result[14]), .C (n_503), .Y (n_510));
  AND2X1 g12602(.A (n_504), .B (query[28]), .Y (n_508));
  AND2X1 g12603(.A (result[14]), .B (n_486), .Y (n_509));
  INVX1 g12604(.A (n_506), .Y (n_507));
  AND2X1 g12605(.A (result[14]), .B (result[15]), .Y (n_506));
  AND2X1 g12606(.A (n_504), .B (n_497), .Y (n_505));
  INVX1 g12607(.A (result[14]), .Y (n_504));
  OAI21X1 g12608(.A (query[30]), .B (n_496), .C (n_503), .Y
       (result[14]));
  OAI21X1 g12609(.A (query[30]), .B (1'b0), .C (query[31]), .Y (n_503));
  OR2X1 g12610(.A (n_497), .B (query[30]), .Y (n_502));
  NOR2X1 g12611(.A (query[27]), .B (query[28]), .Y (n_499));
  OR2X1 g12612(.A (query[15]), .B (query[14]), .Y (n_501));
  OR2X1 g12613(.A (query[25]), .B (query[24]), .Y (n_500));
  INVX1 g12614(.A (result[15]), .Y (n_497));
  AND2X1 g12615(.A (n_486), .B (n_491), .Y (n_496));
  NOR2X1 g12616(.A (query[12]), .B (query[13]), .Y (n_498));
  OR2X1 g12617(.A (query[31]), .B (query[30]), .Y (result[15]));
  INVX1 g12618(.A (query[19]), .Y (n_495));
  INVX1 g12619(.A (query[21]), .Y (n_494));
  INVX1 g12620(.A (query[14]), .Y (n_493));
  INVX1 g12621(.A (query[17]), .Y (n_492));
  INVX1 g12622(.A (query[29]), .Y (n_491));
  INVX1 g12623(.A (query[26]), .Y (n_490));
  INVX1 g12624(.A (query[20]), .Y (n_489));
  INVX1 g12625(.A (query[22]), .Y (n_488));
  INVX1 g12626(.A (query[15]), .Y (n_487));
  INVX1 g12627(.A (query[28]), .Y (n_486));
  INVX1 g12628(.A (query[16]), .Y (n_485));
  INVX1 drc_bufs12654(.A (n_463), .Y (n_470));
  INVX1 drc_bufs12658(.A (n_462), .Y (n_476));
  BUFX2 drc_bufs12664(.A (n_654), .Y (n_460));
  INVX1 drc_bufs12667(.A (n_459), .Y (n_473));
  INVX1 drc_bufs12671(.A (n_458), .Y (n_484));
  INVX1 drc_bufs12683(.A (n_455), .Y (n_478));
  BUFX2 drc_bufs12685(.A (n_752), .Y (n_454));
  BUFX2 drc_bufs12686(.A (n_725), .Y (n_453));
  BUFX2 drc_bufs12687(.A (n_568), .Y (n_452));
  BUFX2 drc_bufs12688(.A (n_499), .Y (n_451));
  BUFX2 drc_bufs12689(.A (n_846), .Y (n_450));
  BUFX2 drc_bufs12690(.A (n_899), .Y (n_449));
  BUFX2 drc_bufs12691(.A (n_555), .Y (n_448));
  BUFX2 drc_bufs12692(.A (n_827), .Y (n_447));
  BUFX2 drc_bufs12693(.A (n_512), .Y (n_446));
  BUFX2 drc_bufs12694(.A (n_633), .Y (n_445));
  BUFX2 drc_bufs12695(.A (n_871), .Y (n_444));
  BUFX2 drc_bufs12696(.A (n_531), .Y (n_443));
  BUFX2 drc_bufs12697(.A (n_874), .Y (n_442));
  BUFX2 drc_bufs12698(.A (n_676), .Y (n_441));
  BUFX2 drc_bufs12699(.A (n_648), .Y (n_440));
  BUFX2 drc_bufs12700(.A (n_848), .Y (n_439));
  BUFX2 drc_bufs12701(.A (n_735), .Y (n_438));
  BUFX2 drc_bufs12702(.A (n_828), .Y (n_437));
  BUFX2 drc_bufs12703(.A (n_577), .Y (n_436));
  BUFX2 drc_bufs12704(.A (n_526), .Y (n_435));
  BUFX2 drc_bufs12705(.A (n_804), .Y (n_434));
  BUFX2 drc_bufs12706(.A (n_895), .Y (n_433));
  BUFX2 drc_bufs12707(.A (n_870), .Y (n_432));
  BUFX2 drc_bufs12708(.A (n_815), .Y (n_431));
  BUFX2 drc_bufs12709(.A (n_789), .Y (n_430));
  BUFX2 drc_bufs12710(.A (n_840), .Y (n_429));
  BUFX2 drc_bufs12711(.A (n_734), .Y (n_428));
  BUFX2 drc_bufs12712(.A (n_522), .Y (n_427));
  BUFX2 drc_bufs12713(.A (n_879), .Y (n_426));
  BUFX2 drc_bufs12714(.A (n_875), .Y (n_425));
  BUFX2 drc_bufs12715(.A (n_683), .Y (n_424));
  BUFX2 drc_bufs12716(.A (n_722), .Y (n_423));
  BUFX2 drc_bufs12717(.A (n_839), .Y (n_422));
  BUFX2 drc_bufs12718(.A (n_803), .Y (n_421));
  BUFX2 drc_bufs12719(.A (n_612), .Y (n_420));
  BUFX2 drc_bufs12720(.A (n_795), .Y (n_419));
  BUFX2 drc_bufs12721(.A (n_533), .Y (n_418));
  BUFX2 drc_bufs12722(.A (n_889), .Y (n_417));
  BUFX2 drc_bufs12723(.A (n_600), .Y (n_416));
  BUFX2 drc_bufs12724(.A (n_556), .Y (n_415));
  BUFX2 drc_bufs12725(.A (n_746), .Y (n_414));
  BUFX2 drc_bufs12726(.A (n_881), .Y (n_413));
  BUFX2 drc_bufs12727(.A (n_702), .Y (n_412));
  BUFX2 drc_bufs12728(.A (n_690), .Y (n_411));
  BUFX2 drc_bufs12729(.A (n_541), .Y (n_410));
  BUFX2 drc_bufs12730(.A (n_751), .Y (n_409));
  BUFX2 drc_bufs12731(.A (n_897), .Y (n_408));
  BUFX2 drc_bufs12732(.A (n_901), .Y (n_407));
  BUFX2 drc_bufs12733(.A (n_628), .Y (n_406));
  BUFX2 drc_bufs12734(.A (n_678), .Y (n_405));
  BUFX2 drc_bufs12735(.A (n_890), .Y (n_404));
  BUFX2 drc_bufs12736(.A (n_675), .Y (n_403));
  BUFX2 drc_bufs12737(.A (n_629), .Y (n_402));
  BUFX2 drc_bufs12738(.A (n_635), .Y (n_401));
  BUFX2 drc_bufs12739(.A (n_517), .Y (n_400));
  BUFX2 drc_bufs12740(.A (n_750), .Y (n_399));
  BUFX2 drc_bufs12741(.A (n_688), .Y (n_398));
  BUFX2 drc_bufs12742(.A (n_764), .Y (n_397));
  BUFX2 drc_bufs12743(.A (n_670), .Y (n_396));
  BUFX2 drc_bufs12744(.A (n_816), .Y (n_395));
  BUFX2 drc_bufs12745(.A (n_544), .Y (n_394));
  BUFX2 drc_bufs12746(.A (n_666), .Y (n_393));
  BUFX2 drc_bufs12747(.A (n_894), .Y (n_458));
  BUFX2 drc_bufs12748(.A (n_713), .Y (n_461));
  BUFX2 drc_bufs12749(.A (n_699), .Y (n_455));
  BUFX2 drc_bufs12750(.A (n_551), .Y (n_464));
  BUFX2 drc_bufs12751(.A (n_529), .Y (n_468));
  BUFX2 drc_bufs12752(.A (n_516), .Y (n_463));
  BUFX2 drc_bufs12753(.A (n_498), .Y (n_466));
  BUFX2 drc_bufs12754(.A (n_677), .Y (n_462));
  BUFX2 drc_bufs12755(.A (n_650), .Y (n_457));
  BUFX2 drc_bufs12756(.A (n_647), .Y (n_467));
  BUFX2 drc_bufs12757(.A (n_615), .Y (n_469));
  BUFX2 drc_bufs12758(.A (n_597), .Y (n_459));
  BUFX2 drc_bufs12759(.A (n_576), .Y (n_465));
  BUFX2 drc_bufs12760(.A (n_557), .Y (n_456));
  XOR2X1 g2(.A (n_845), .B (n_821), .Y (n_392));
  XOR2X1 g12838(.A (n_655), .B (n_651), .Y (n_391));
  AND2X1 g3070(.A (result[4]), .B (result[14]), .Y
       (\genblk1[12].inst_n_710 ));
  AND2X1 g3071(.A (result[4]), .B (result[15]), .Y
       (\genblk1[12].inst_n_709 ));
  AND2X1 g3072(.A (result[4]), .B (n_346), .Y (\genblk1[12].inst_n_713
       ));
  AND2X1 g3073(.A (result[4]), .B (result[13]), .Y
       (\genblk1[12].inst_n_711 ));
  AND2X1 g3074(.A (result[4]), .B (result[12]), .Y
       (\genblk1[12].inst_n_712 ));
  AND2X1 g3075(.A (result[4]), .B (result[10]), .Y
       (\genblk1[12].inst_n_714 ));
  AND2X1 g3076(.A (result[4]), .B (result[9]), .Y
       (\genblk1[12].inst_n_715 ));
  AND2X1 g3077(.A (result[4]), .B (result[8]), .Y
       (\genblk1[12].inst_n_716 ));
  AND2X1 g3078(.A (result[4]), .B (result[7]), .Y
       (\genblk1[12].inst_n_717 ));
  AND2X1 g3079(.A (result[4]), .B (result[6]), .Y
       (\genblk1[12].inst_n_718 ));
  AND2X1 g3080(.A (result[4]), .B (result[5]), .Y
       (\genblk1[12].inst_n_719 ));
  OR2X1 g3081(.A (n_390), .B (n_365), .Y (result[4]));
  OR2X1 g3082(.A (n_329), .B (n_376), .Y (n_390));
  NAND3X1 g3083(.A (n_330), .B (n_343), .C (n_334), .Y (n_389));
  AOI22X1 g3084(.A (n_387), .B (n_361), .C (n_344), .D (\eps[11] [20]),
       .Y (n_388));
  NOR3X1 g3085(.A (n_386), .B (n_339), .C (n_366), .Y (n_387));
  OAI21X1 g3086(.A (\genblk1[15].inst_n_1114 ), .B (\eps[11] [16]), .C
       (n_324), .Y (n_386));
  AOI21X1 g3087(.A (result[10]), .B (n_331), .C (n_326), .Y (n_385));
  NAND2X1 g3088(.A (\eps[11] [15]), .B (n_338), .Y (n_384));
  NOR2X1 g3089(.A (\eps[11] [15]), .B (n_338), .Y (n_383));
  AOI21X1 g3090(.A (result[9]), .B (n_352), .C (n_328), .Y (n_382));
  AOI21X1 g3091(.A (n_348), .B (\eps[11] [14]), .C (n_380), .Y (n_381));
  OAI21X1 g3092(.A (result[8]), .B (n_378), .C (n_379), .Y (n_380));
  OAI21X1 g3093(.A (n_357), .B (n_377), .C (\eps[11] [13]), .Y (n_379));
  NOR3X1 g3094(.A (n_357), .B (\eps[11] [13]), .C (n_377), .Y (n_378));
  AND2X1 g3095(.A (n_325), .B (n_358), .Y (n_377));
  OAI21X1 g3096(.A (result[14]), .B (n_368), .C (n_374), .Y (n_376));
  AOI21X1 g3097(.A (result[6]), .B (n_332), .C (n_327), .Y (n_375));
  OAI21X1 g3098(.A (n_369), .B (n_370), .C (n_336), .Y (n_374));
  NOR2X1 g3099(.A (\eps[11] [11]), .B (n_337), .Y (n_373));
  NAND2X1 g3100(.A (\eps[11] [11]), .B (n_337), .Y (n_372));
  AOI22X1 g3101(.A (n_333), .B (n_353), .C (result[5]), .D (n_349), .Y
       (n_371));
  NOR3X1 g3102(.A (n_360), .B (n_335), .C (n_366), .Y (n_370));
  NOR3X1 g3103(.A (result[13]), .B (n_351), .C (n_359), .Y (n_369));
  OR2X1 g3104(.A (n_359), .B (n_350), .Y (n_368));
  AOI21X1 g3105(.A (n_345), .B (\eps[11] [10]), .C (query[9]), .Y
       (n_367));
  INVX1 g3106(.A (n_323), .Y (n_366));
  OR2X1 g3107(.A (n_355), .B (n_354), .Y (n_365));
  AOI22X1 g3108(.A (\eps[11] [17]), .B (n_340), .C
       (\genblk1[15].inst_n_1114 ), .D (\eps[11] [16]), .Y (n_364));
  AOI21X1 g3109(.A (result[13]), .B (n_351), .C (n_359), .Y (n_363));
  INVX1 g3111(.A (n_360), .Y (n_361));
  OR2X1 g3112(.A (\eps[11] [12]), .B (n_347), .Y (n_358));
  NAND2X1 g3113(.A (result[14]), .B (n_350), .Y (n_362));
  AND2X1 g3114(.A (n_341), .B (result[12]), .Y (n_360));
  AND2X1 g3115(.A (n_342), .B (result[15]), .Y (n_359));
  NOR2X1 g3116(.A (1'b0), .B (1'b0), .Y (n_356));
  OR2X1 g3117(.A (1'b0), .B (1'b0), .Y (n_355));
  OR2X1 g3118(.A (1'b0), .B (\eps[11] [21]), .Y (n_354));
  AND2X1 g3119(.A (\eps[11] [12]), .B (n_347), .Y (n_357));
  INVX1 g3120(.A (query[8]), .Y (n_353));
  INVX1 g3121(.A (\eps[11] [14]), .Y (n_352));
  INVX1 g3122(.A (\eps[11] [18]), .Y (n_351));
  INVX1 g3123(.A (\eps[11] [19]), .Y (n_350));
  INVX1 g3124(.A (\eps[11] [10]), .Y (n_349));
  INVX1 g3125(.A (result[9]), .Y (n_348));
  INVX1 g3126(.A (result[7]), .Y (n_347));
  INVX1 g3127(.A (\genblk1[15].inst_n_1114 ), .Y (n_346));
  INVX1 g3128(.A (result[5]), .Y (n_345));
  INVX1 g3129(.A (result[15]), .Y (n_344));
  INVX1 g3130(.A (\eps[11] [31]), .Y (n_343));
  INVX1 g3131(.A (\eps[11] [20]), .Y (n_342));
  INVX1 g3132(.A (\eps[11] [17]), .Y (n_341));
  INVX1 g3133(.A (result[12]), .Y (n_340));
  INVX1 drc_bufs3143(.A (n_336), .Y (n_339));
  BUFX2 drc_bufs3145(.A (n_364), .Y (n_335));
  BUFX2 drc_bufs3146(.A (n_356), .Y (n_334));
  BUFX2 drc_bufs3147(.A (n_367), .Y (n_333));
  BUFX2 drc_bufs3148(.A (n_372), .Y (n_332));
  BUFX2 drc_bufs3149(.A (n_384), .Y (n_331));
  BUFX2 drc_bufs3150(.A (n_388), .Y (n_330));
  BUFX2 drc_bufs3151(.A (n_389), .Y (n_329));
  BUFX2 drc_bufs3152(.A (n_381), .Y (n_328));
  BUFX2 drc_bufs3153(.A (n_373), .Y (n_327));
  BUFX2 drc_bufs3154(.A (n_383), .Y (n_326));
  BUFX2 drc_bufs3155(.A (n_375), .Y (n_325));
  BUFX2 drc_bufs3156(.A (n_385), .Y (n_324));
  BUFX2 drc_bufs3157(.A (n_363), .Y (n_323));
  BUFX2 drc_bufs3158(.A (n_382), .Y (n_338));
  BUFX2 drc_bufs3159(.A (n_371), .Y (n_337));
  BUFX2 drc_bufs3160(.A (n_362), .Y (n_336));
  AND2X1 g3141(.A (result[5]), .B (result[13]), .Y
       (\genblk1[11].inst_n_710 ));
  AND2X1 g3142(.A (result[5]), .B (result[15]), .Y
       (\genblk1[11].inst_n_708 ));
  AND2X1 g3143(.A (result[5]), .B (n_275), .Y (\genblk1[11].inst_n_712
       ));
  AND2X1 g3144(.A (result[5]), .B (result[12]), .Y
       (\genblk1[11].inst_n_711 ));
  AND2X1 g3145(.A (result[5]), .B (result[14]), .Y
       (\genblk1[11].inst_n_709 ));
  AND2X1 g3146(.A (result[5]), .B (result[8]), .Y
       (\genblk1[11].inst_n_715 ));
  AND2X1 g3147(.A (result[5]), .B (result[9]), .Y
       (\genblk1[11].inst_n_714 ));
  AND2X1 g3148(.A (result[5]), .B (result[10]), .Y
       (\genblk1[11].inst_n_713 ));
  AND2X1 g3149(.A (result[5]), .B (result[7]), .Y
       (\genblk1[11].inst_n_716 ));
  AND2X1 g3150(.A (result[5]), .B (result[6]), .Y
       (\genblk1[11].inst_n_717 ));
  OR2X1 g3151(.A (n_268), .B (n_309), .Y (result[5]));
  NAND3X1 g3152(.A (n_281), .B (n_270), .C (n_318), .Y (n_322));
  NAND3X1 g3153(.A (n_320), .B (n_298), .C (n_307), .Y (n_321));
  OAI21X1 g3154(.A (result[8]), .B (n_269), .C (n_262), .Y (n_320));
  AOI22X1 g3155(.A (n_317), .B (n_291), .C (n_283), .D (\eps[10] [15]),
       .Y (n_319));
  NOR3X1 g3156(.A (n_316), .B (1'b0), .C (n_313), .Y (n_318));
  AND2X1 g3157(.A (n_263), .B (n_289), .Y (n_317));
  OR2X1 g3158(.A (n_314), .B (1'b0), .Y (n_316));
  AOI21X1 g3159(.A (result[8]), .B (n_280), .C (n_264), .Y (n_315));
  AND2X1 g3160(.A (n_300), .B (n_310), .Y (n_314));
  AND2X1 g3161(.A (n_307), .B (n_308), .Y (n_313));
  AOI21X1 g3162(.A (n_277), .B (\eps[10] [13]), .C (n_265), .Y (n_312));
  AOI22X1 g3163(.A (n_271), .B (n_282), .C (result[6]), .D (n_279), .Y
       (n_311));
  OAI21X1 g3164(.A (result[13]), .B (n_286), .C (n_305), .Y (n_310));
  OAI21X1 g3165(.A (result[15]), .B (n_287), .C (n_306), .Y (n_309));
  OAI21X1 g3166(.A (result[10]), .B (n_272), .C (n_261), .Y (n_308));
  AND2X1 g3167(.A (n_300), .B (n_299), .Y (n_307));
  OR2X1 g3168(.A (n_267), .B (result[14]), .Y (n_306));
  OR2X1 g3169(.A (n_266), .B (result[12]), .Y (n_305));
  NAND2X1 g3170(.A (\eps[10] [14]), .B (n_291), .Y (n_304));
  NAND2X1 g3171(.A (\eps[10] [16]), .B (n_292), .Y (n_303));
  NAND2X1 g3172(.A (\eps[10] [20]), .B (n_274), .Y (n_302));
  NAND2X1 g3173(.A (\eps[10] [18]), .B (n_273), .Y (n_301));
  AND2X1 g3174(.A (n_273), .B (n_295), .Y (n_299));
  AND2X1 g3175(.A (n_292), .B (n_293), .Y (n_298));
  AOI21X1 g3176(.A (n_285), .B (\eps[10] [12]), .C (query[11]), .Y
       (n_297));
  AND2X1 g3177(.A (n_274), .B (n_294), .Y (n_300));
  OR2X1 g3178(.A (\eps[10] [18]), .B (n_284), .Y (n_295));
  OR2X1 g3179(.A (\eps[10] [20]), .B (n_278), .Y (n_294));
  OR2X1 g3180(.A (\eps[10] [16]), .B (n_276), .Y (n_293));
  NAND2X1 g3181(.A (result[15]), .B (n_287), .Y (n_296));
  OR2X1 g3182(.A (\eps[10] [13]), .B (n_277), .Y (n_289));
  NAND2X1 g3183(.A (\genblk1[15].inst_n_1114 ), .B (\eps[10] [17]), .Y
       (n_288));
  OR2X1 g3184(.A (\eps[10] [17]), .B (\genblk1[15].inst_n_1114 ), .Y
       (n_292));
  OR2X1 g3185(.A (\eps[10] [15]), .B (n_283), .Y (n_291));
  NAND2X1 g3186(.A (result[13]), .B (n_286), .Y (n_290));
  INVX1 g3187(.A (\eps[10] [21]), .Y (n_287));
  INVX1 g3188(.A (\eps[10] [19]), .Y (n_286));
  INVX1 g3189(.A (result[6]), .Y (n_285));
  INVX1 g3190(.A (result[12]), .Y (n_284));
  INVX1 g3191(.A (result[9]), .Y (n_283));
  INVX1 g3192(.A (query[10]), .Y (n_282));
  INVX1 g3193(.A (\eps[10] [22]), .Y (n_281));
  INVX1 g3194(.A (\eps[10] [14]), .Y (n_280));
  INVX1 g3195(.A (\eps[10] [12]), .Y (n_279));
  INVX1 g3196(.A (result[14]), .Y (n_278));
  INVX1 g3197(.A (result[7]), .Y (n_277));
  INVX1 g3198(.A (result[10]), .Y (n_276));
  INVX1 g3199(.A (\genblk1[15].inst_n_1114 ), .Y (n_275));
  BUFX2 drc_bufs3207(.A (n_303), .Y (n_272));
  BUFX2 drc_bufs3208(.A (n_297), .Y (n_271));
  BUFX2 drc_bufs3209(.A (n_321), .Y (n_270));
  BUFX2 drc_bufs3210(.A (n_304), .Y (n_269));
  BUFX2 drc_bufs3211(.A (n_322), .Y (n_268));
  BUFX2 drc_bufs3212(.A (n_302), .Y (n_267));
  BUFX2 drc_bufs3213(.A (n_301), .Y (n_266));
  BUFX2 drc_bufs3214(.A (n_311), .Y (n_265));
  BUFX2 drc_bufs3215(.A (n_312), .Y (n_264));
  BUFX2 drc_bufs3216(.A (n_315), .Y (n_263));
  BUFX2 drc_bufs3217(.A (n_319), .Y (n_262));
  BUFX2 drc_bufs3218(.A (n_288), .Y (n_261));
  BUFX2 drc_bufs3219(.A (n_296), .Y (n_274));
  BUFX2 drc_bufs3220(.A (n_290), .Y (n_273));
  NAND3X1 g3476(.A (n_222), .B (n_186), .C (n_260), .Y (result[0]));
  NOR3X1 g3477(.A (1'b0), .B (\eps[15] [29]), .C (n_189), .Y (n_260));
  NAND3X1 g3478(.A (n_183), .B (n_224), .C (n_218), .Y (n_259));
  AOI21X1 g3479(.A (n_215), .B (n_257), .C (1'b0), .Y (n_258));
  OAI21X1 g3480(.A (n_256), .B (n_230), .C (n_244), .Y (n_257));
  OAI21X1 g3481(.A (\genblk1[15].inst_n_1114 ), .B (\eps[15] [12]), .C
       (n_255), .Y (n_256));
  OAI21X1 g3482(.A (result[9]), .B (n_188), .C (n_174), .Y (n_255));
  AOI22X1 g3483(.A (n_253), .B (n_221), .C (n_201), .D (\eps[15] [11]),
       .Y (n_254));
  OAI21X1 g3484(.A (result[8]), .B (n_195), .C (n_252), .Y (n_253));
  INVX1 g3485(.A (n_171), .Y (n_252));
  AOI21X1 g3486(.A (result[8]), .B (n_195), .C (n_180), .Y (n_251));
  AOI21X1 g3487(.A (\eps[15] [8]), .B (n_184), .C (n_177), .Y (n_250));
  AOI21X1 g3488(.A (n_247), .B (n_246), .C (result[7]), .Y (n_249));
  NAND3X1 g3489(.A (n_247), .B (n_241), .C (n_190), .Y (n_248));
  OR2X1 g3490(.A (n_231), .B (n_245), .Y (n_247));
  NOR3X1 g3491(.A (\eps[15] [8]), .B (n_240), .C (n_191), .Y (n_246));
  OAI21X1 g3492(.A (n_198), .B (\eps[15] [4]), .C (n_172), .Y (n_245));
  AND2X1 g3493(.A (n_176), .B (n_233), .Y (n_244));
  AOI21X1 g3495(.A (result[2]), .B (n_204), .C (n_181), .Y (n_242));
  AOI22X1 g3496(.A (n_236), .B (n_198), .C (n_192), .D (\eps[15] [7]),
       .Y (n_243));
  INVX1 g3497(.A (n_240), .Y (n_241));
  OAI21X1 g3498(.A (result[4]), .B (n_185), .C (n_229), .Y (n_240));
  AOI21X1 g3499(.A (n_208), .B (\eps[15] [3]), .C (n_179), .Y (n_239));
  AOI21X1 g3500(.A (n_202), .B (\eps[15] [15]), .C (n_178), .Y (n_238));
  NOR2X1 g3501(.A (n_175), .B (n_230), .Y (n_237));
  AND2X1 g3502(.A (n_232), .B (\eps[15] [4]), .Y (n_236));
  AOI22X1 g3503(.A (n_187), .B (n_200), .C (result[1]), .D (n_207), .Y
       (n_235));
  NAND2X1 g3504(.A (\eps[15] [5]), .B (n_223), .Y (n_234));
  OR2X1 g3505(.A (n_228), .B (result[13]), .Y (n_233));
  INVX1 g3506(.A (n_231), .Y (n_232));
  OR2X1 g3507(.A (n_182), .B (result[5]), .Y (n_229));
  OAI21X1 g3508(.A (n_206), .B (\eps[15] [5]), .C (n_223), .Y (n_231));
  OAI21X1 g3509(.A (n_202), .B (\eps[15] [15]), .C (n_173), .Y (n_230));
  OAI21X1 g3510(.A (n_202), .B (\eps[15] [15]), .C (\eps[15] [14]), .Y
       (n_228));
  NAND2X1 g3511(.A (\eps[15] [6]), .B (n_213), .Y (n_227));
  NAND2X1 g3512(.A (\eps[15] [10]), .B (n_217), .Y (n_226));
  AOI21X1 g3513(.A (n_194), .B (\eps[15] [2]), .C (query[1]), .Y
       (n_225));
  NOR3X1 g3514(.A (n_210), .B (\eps[15] [25]), .C (\eps[15] [26]), .Y
       (n_224));
  NOR3X1 g3515(.A (n_212), .B (\eps[15] [19]), .C (\eps[15] [20]), .Y
       (n_222));
  AND2X1 g3516(.A (n_217), .B (n_216), .Y (n_221));
  AOI22X1 g3517(.A (n_197), .B (result[12]), .C (result[13]), .D
       (n_203), .Y (n_220));
  AOI22X1 g12839(.A (\eps[15] [13]), .B (n_196), .C
       (\genblk1[15].inst_n_1114 ), .D (\eps[15] [12]), .Y (n_219));
  NOR3X1 g12840(.A (n_214), .B (1'b0), .C (\eps[15] [28]), .Y (n_218));
  AND2X1 g12841(.A (n_213), .B (n_211), .Y (n_223));
  OR2X1 g12842(.A (\eps[15] [10]), .B (n_205), .Y (n_216));
  OR2X1 g12843(.A (\eps[15] [16]), .B (n_199), .Y (n_215));
  AND2X1 g12844(.A (\eps[15] [16]), .B (n_199), .Y (n_214));
  OR2X1 g12845(.A (\eps[15] [11]), .B (n_201), .Y (n_217));
  OR2X1 g12846(.A (\eps[15] [18]), .B (\eps[15] [17]), .Y (n_212));
  OR2X1 g12847(.A (\eps[15] [6]), .B (n_193), .Y (n_211));
  OR2X1 g12848(.A (1'b0), .B (\eps[15] [23]), .Y (n_210));
  NOR2X1 g12849(.A (\eps[15] [31]), .B (1'b0), .Y (n_209));
  OR2X1 g12850(.A (\eps[15] [7]), .B (n_192), .Y (n_213));
  INVX1 g12851(.A (result[2]), .Y (n_208));
  INVX1 g12852(.A (\eps[15] [2]), .Y (n_207));
  INVX1 g12853(.A (result[4]), .Y (n_206));
  INVX1 g12854(.A (result[9]), .Y (n_205));
  INVX1 g12855(.A (\eps[15] [3]), .Y (n_204));
  INVX1 g12856(.A (\eps[15] [14]), .Y (n_203));
  INVX1 g12857(.A (result[14]), .Y (n_202));
  INVX1 g12858(.A (result[10]), .Y (n_201));
  INVX1 g12859(.A (\genblk1[15].inst_n_1114 ), .Y (result[11]));
  INVX1 g12860(.A (query[0]), .Y (n_200));
  INVX1 g12861(.A (result[15]), .Y (n_199));
  INVX1 g12862(.A (result[3]), .Y (n_198));
  INVX1 g12863(.A (\eps[15] [13]), .Y (n_197));
  INVX1 g12864(.A (result[12]), .Y (n_196));
  INVX1 g12865(.A (\eps[15] [9]), .Y (n_195));
  INVX1 g12866(.A (result[1]), .Y (n_194));
  INVX1 g12867(.A (result[5]), .Y (n_193));
  INVX1 g12868(.A (result[6]), .Y (n_192));
  INVX1 drc_bufs3549(.A (n_190), .Y (n_191));
  BUFX2 drc_bufs3551(.A (n_259), .Y (n_189));
  BUFX2 drc_bufs3552(.A (n_226), .Y (n_188));
  BUFX2 drc_bufs3553(.A (n_225), .Y (n_187));
  BUFX2 drc_bufs3554(.A (n_209), .Y (n_186));
  BUFX2 drc_bufs3555(.A (n_234), .Y (n_185));
  BUFX2 drc_bufs3556(.A (n_248), .Y (n_184));
  BUFX2 drc_bufs3557(.A (n_258), .Y (n_183));
  BUFX2 drc_bufs3558(.A (n_227), .Y (n_182));
  BUFX2 drc_bufs3559(.A (n_239), .Y (n_181));
  BUFX2 drc_bufs3560(.A (n_250), .Y (n_180));
  BUFX2 drc_bufs3561(.A (n_235), .Y (n_179));
  BUFX2 drc_bufs3562(.A (n_237), .Y (n_178));
  BUFX2 drc_bufs3563(.A (n_249), .Y (n_177));
  BUFX2 drc_bufs3564(.A (n_238), .Y (n_176));
  BUFX2 drc_bufs3565(.A (n_219), .Y (n_175));
  BUFX2 drc_bufs3566(.A (n_254), .Y (n_174));
  BUFX2 drc_bufs3567(.A (n_220), .Y (n_173));
  BUFX2 drc_bufs3568(.A (n_242), .Y (n_172));
  BUFX2 drc_bufs3569(.A (n_251), .Y (n_171));
  BUFX2 drc_bufs3570(.A (n_243), .Y (n_190));
  NOR2X1 g12869(.A (\genblk1[15].inst_n_1114 ), .B (n_169), .Y (n_170));
  AND2X1 g12870(.A (result[3]), .B (result[15]), .Y
       (\genblk1[13].inst_n_710 ));
  AND2X1 g12871(.A (result[3]), .B (result[14]), .Y
       (\genblk1[13].inst_n_711 ));
  AND2X1 g12872(.A (result[3]), .B (result[13]), .Y
       (\genblk1[13].inst_n_712 ));
  AND2X1 g12873(.A (result[3]), .B (result[6]), .Y
       (\genblk1[13].inst_n_719 ));
  AND2X1 g12874(.A (result[3]), .B (result[12]), .Y
       (\genblk1[13].inst_n_713 ));
  AND2X1 g12875(.A (result[3]), .B (result[10]), .Y
       (\genblk1[13].inst_n_715 ));
  AND2X1 g12876(.A (result[3]), .B (result[9]), .Y
       (\genblk1[13].inst_n_716 ));
  AND2X1 g12877(.A (result[3]), .B (result[8]), .Y
       (\genblk1[13].inst_n_717 ));
  AND2X1 g12878(.A (result[3]), .B (result[7]), .Y
       (\genblk1[13].inst_n_718 ));
  AND2X1 g12879(.A (result[3]), .B (result[5]), .Y
       (\genblk1[13].inst_n_720 ));
  AND2X1 g12880(.A (result[3]), .B (result[4]), .Y
       (\genblk1[13].inst_n_721 ));
  INVX1 g12881(.A (result[3]), .Y (n_169));
  OR2X1 g12882(.A (n_101), .B (n_95), .Y (result[3]));
  NAND3X1 g12883(.A (n_136), .B (n_104), .C (n_167), .Y (n_168));
  AND2X1 g12884(.A (n_116), .B (n_93), .Y (n_167));
  NAND3X1 g12885(.A (n_127), .B (n_133), .C (n_106), .Y (n_166));
  AOI21X1 g12886(.A (result[14]), .B (n_115), .C (n_94), .Y (n_165));
  AOI21X1 g12887(.A (n_121), .B (\eps[12] [17]), .C (n_96), .Y (n_164));
  AOI22X1 g12888(.A (n_162), .B (n_103), .C (result[12]), .D (n_114),
       .Y (n_163));
  NOR3X1 g12889(.A (n_151), .B (n_107), .C (n_161), .Y (n_162));
  OAI21X1 g12890(.A (n_149), .B (n_139), .C (n_160), .Y (n_161));
  OAI21X1 g12891(.A (query[6]), .B (query[7]), .C (n_157), .Y (n_160));
  AOI22X1 g12892(.A (n_155), .B (\eps[12] [8]), .C (n_119), .D
       (\eps[12] [16]), .Y (n_159));
  AOI21X1 g12893(.A (n_150), .B (n_152), .C (n_146), .Y (n_158));
  INVX1 g12894(.A (n_91), .Y (n_157));
  AOI21X1 g12895(.A (\eps[12] [8]), .B (n_153), .C (n_155), .Y (n_156));
  AND2X1 g12896(.A (n_153), .B (n_122), .Y (n_155));
  NAND3X1 g12897(.A (n_99), .B (n_147), .C (n_105), .Y (n_154));
  OR2X1 g12898(.A (n_148), .B (result[5]), .Y (n_152));
  NOR3X1 g12899(.A (n_130), .B (n_138), .C (n_146), .Y (n_153));
  OAI21X1 g12900(.A (result[10]), .B (n_102), .C (n_92), .Y (n_151));
  AND2X1 g12901(.A (n_145), .B (n_132), .Y (n_150));
  AND2X1 g12902(.A (n_144), .B (n_131), .Y (n_149));
  OR2X1 g12903(.A (n_138), .B (n_113), .Y (n_148));
  OR2X1 g12904(.A (n_97), .B (result[14]), .Y (n_147));
  OR2X1 g12905(.A (n_100), .B (result[6]), .Y (n_145));
  OR2X1 g12906(.A (n_98), .B (result[8]), .Y (n_144));
  OR2X1 g12907(.A (n_139), .B (n_137), .Y (n_146));
  NAND2X1 g12908(.A (\eps[12] [10]), .B (n_134), .Y (n_143));
  NAND2X1 g12909(.A (\eps[12] [12]), .B (n_135), .Y (n_142));
  NAND2X1 g12910(.A (\eps[12] [14]), .B (n_129), .Y (n_141));
  NAND2X1 g12911(.A (\eps[12] [18]), .B (n_133), .Y (n_140));
  OAI21X1 g12912(.A (n_108), .B (\eps[12] [12]), .C (n_135), .Y
       (n_137));
  NOR3X1 g12913(.A (1'b0), .B (1'b0), .C (n_128), .Y (n_136));
  OAI21X1 g12914(.A (n_120), .B (\eps[12] [14]), .C (n_129), .Y
       (n_139));
  OAI21X1 g12915(.A (n_109), .B (\eps[12] [10]), .C (n_134), .Y
       (n_138));
  OR2X1 g12916(.A (n_111), .B (result[7]), .Y (n_132));
  OR2X1 g12917(.A (n_112), .B (result[9]), .Y (n_131));
  AND2X1 g12918(.A (n_113), .B (result[5]), .Y (n_130));
  OR2X1 g12919(.A (\eps[12] [13]), .B (n_117), .Y (n_135));
  OR2X1 g12920(.A (\eps[12] [11]), .B (n_110), .Y (n_134));
  OR2X1 g12921(.A (\eps[12] [19]), .B (n_118), .Y (n_133));
  OR2X1 g12922(.A (1'b0), .B (1'b0), .Y (n_128));
  OR2X1 g3200(.A (\eps[12] [17]), .B (n_121), .Y (n_127));
  NAND2X1 g3201(.A (n_118), .B (\eps[12] [19]), .Y (n_126));
  NAND2X1 g3202(.A (\genblk1[15].inst_n_1114 ), .B (\eps[12] [15]), .Y
       (n_125));
  NOR2X1 g3203(.A (\eps[12] [20]), .B (1'b0), .Y (n_124));
  NOR2X1 g3204(.A (1'b0), .B (1'b0), .Y (n_123));
  OR2X1 g3205(.A (\eps[12] [15]), .B (\genblk1[15].inst_n_1114 ), .Y
       (n_129));
  INVX1 g3206(.A (result[4]), .Y (n_122));
  INVX1 g3207(.A (result[13]), .Y (n_121));
  INVX1 g3208(.A (result[10]), .Y (n_120));
  INVX1 g3209(.A (result[12]), .Y (n_119));
  INVX1 g3210(.A (result[15]), .Y (n_118));
  INVX1 g3211(.A (result[9]), .Y (n_117));
  INVX1 g3212(.A (\eps[12] [31]), .Y (n_116));
  INVX1 g3213(.A (\eps[12] [18]), .Y (n_115));
  INVX1 g3214(.A (\eps[12] [16]), .Y (n_114));
  INVX1 g3215(.A (\eps[12] [9]), .Y (n_113));
  INVX1 g3216(.A (\eps[12] [13]), .Y (n_112));
  INVX1 g3217(.A (\eps[12] [11]), .Y (n_111));
  INVX1 g3218(.A (result[7]), .Y (n_110));
  INVX1 g3219(.A (result[6]), .Y (n_109));
  INVX1 g3220(.A (result[8]), .Y (n_108));
  BUFX2 drc_bufs(.A (n_158), .Y (n_107));
  BUFX2 drc_bufs3221(.A (n_165), .Y (n_106));
  BUFX2 drc_bufs3222(.A (n_124), .Y (n_105));
  BUFX2 drc_bufs3223(.A (n_123), .Y (n_104));
  BUFX2 drc_bufs3224(.A (n_159), .Y (n_103));
  BUFX2 drc_bufs3225(.A (n_141), .Y (n_102));
  BUFX2 drc_bufs3226(.A (n_168), .Y (n_101));
  BUFX2 drc_bufs3227(.A (n_143), .Y (n_100));
  BUFX2 drc_bufs3228(.A (n_126), .Y (n_99));
  BUFX2 drc_bufs3229(.A (n_142), .Y (n_98));
  BUFX2 drc_bufs3230(.A (n_140), .Y (n_97));
  BUFX2 drc_bufs3231(.A (n_163), .Y (n_96));
  BUFX2 drc_bufs3232(.A (n_154), .Y (n_95));
  BUFX2 drc_bufs3233(.A (n_164), .Y (n_94));
  BUFX2 drc_bufs3234(.A (n_166), .Y (n_93));
  BUFX2 drc_bufs3235(.A (n_125), .Y (n_92));
  BUFX2 drc_bufs3236(.A (n_156), .Y (n_91));
  BUFX2 drc_bufs3237(.A (n_170), .Y (\genblk1[13].inst_n_714 ));
  AND2X1 g3446(.A (result[1]), .B (result[5]), .Y
       (\genblk1[15].inst_n_722 ));
  AND2X1 g3447(.A (result[1]), .B (result[9]), .Y
       (\genblk1[15].inst_n_718 ));
  AND2X1 g3448(.A (result[1]), .B (result[2]), .Y
       (\genblk1[15].inst_n_725 ));
  AND2X1 g3449(.A (result[1]), .B (result[8]), .Y
       (\genblk1[15].inst_n_719 ));
  AND2X1 g3450(.A (result[1]), .B (result[7]), .Y
       (\genblk1[15].inst_n_720 ));
  AND2X1 g3451(.A (result[1]), .B (result[6]), .Y
       (\genblk1[15].inst_n_721 ));
  NOR2X1 g3452(.A (\genblk1[15].inst_n_1114 ), .B (n_89), .Y (n_90));
  AND2X1 g3453(.A (result[1]), .B (result[10]), .Y
       (\genblk1[15].inst_n_717 ));
  AND2X1 g3454(.A (result[1]), .B (result[3]), .Y
       (\genblk1[15].inst_n_724 ));
  AND2X1 g3455(.A (result[1]), .B (result[15]), .Y
       (\genblk1[15].inst_n_712 ));
  AND2X1 g3456(.A (result[1]), .B (result[14]), .Y
       (\genblk1[15].inst_n_713 ));
  AND2X1 g3457(.A (result[1]), .B (result[13]), .Y
       (\genblk1[15].inst_n_714 ));
  AND2X1 g3458(.A (result[1]), .B (result[12]), .Y
       (\genblk1[15].inst_n_715 ));
  AND2X1 g3459(.A (result[1]), .B (result[4]), .Y
       (\genblk1[15].inst_n_723 ));
  INVX1 g3460(.A (result[1]), .Y (n_89));
  OR2X1 g3461(.A (n_9), .B (n_7), .Y (result[1]));
  NAND3X1 g3462(.A (n_11), .B (n_15), .C (n_55), .Y (n_88));
  AOI21X1 g3463(.A (n_46), .B (n_86), .C (\eps[14] [18]), .Y (n_87));
  OAI21X1 g3464(.A (result[14]), .B (n_83), .C (n_1), .Y (n_86));
  NAND2X1 g3465(.A (\eps[14] [16]), .B (n_3), .Y (n_85));
  NAND2X1 g3466(.A (result[14]), .B (n_83), .Y (n_84));
  NOR3X1 g3467(.A (n_69), .B (n_20), .C (n_82), .Y (n_83));
  NOR3X1 g3468(.A (n_17), .B (n_81), .C (n_54), .Y (n_82));
  OAI21X1 g3469(.A (n_25), .B (\eps[14] [12]), .C (n_2), .Y (n_81));
  NAND3X1 g3470(.A (n_66), .B (n_71), .C (n_19), .Y (n_80));
  AOI22X1 g3471(.A (n_52), .B (n_16), .C (n_33), .D (\eps[14] [11]), .Y
       (n_79));
  AOI21X1 g3472(.A (result[7]), .B (n_26), .C (n_6), .Y (n_78));
  AOI21X1 g3473(.A (n_30), .B (\eps[14] [8]), .C (n_5), .Y (n_77));
  AOI22X1 g3474(.A (n_75), .B (n_72), .C (result[6]), .D (n_29), .Y
       (n_76));
  NOR3X1 g3475(.A (n_68), .B (n_70), .C (n_73), .Y (n_75));
  AOI21X1 g12923(.A (n_14), .B (n_63), .C (n_54), .Y (n_74));
  NOR3X1 g12924(.A (result[2]), .B (n_27), .C (n_64), .Y (n_73));
  OR2X1 g12925(.A (n_64), .B (n_50), .Y (n_72));
  OR2X1 g12926(.A (n_10), .B (result[7]), .Y (n_71));
  NOR3X1 g12927(.A (result[3]), .B (n_28), .C (n_53), .Y (n_70));
  OAI21X1 g12928(.A (result[13]), .B (n_34), .C (n_61), .Y (n_69));
  OAI21X1 g12929(.A (result[5]), .B (n_35), .C (n_62), .Y (n_68));
  NAND2X1 g12930(.A (\eps[14] [9]), .B (n_52), .Y (n_67));
  OR2X1 g12931(.A (n_13), .B (result[8]), .Y (n_66));
  NAND3X1 g12932(.A (n_47), .B (n_51), .C (n_18), .Y (n_65));
  INVX1 g12933(.A (n_0), .Y (n_64));
  OR2X1 g12934(.A (n_56), .B (result[10]), .Y (n_63));
  OR2X1 g12935(.A (n_8), .B (result[4]), .Y (n_62));
  OR2X1 g12936(.A (n_12), .B (result[12]), .Y (n_61));
  AOI21X1 g12937(.A (result[3]), .B (n_28), .C (n_53), .Y (n_60));
  NAND2X1 g12938(.A (\eps[14] [6]), .B (n_22), .Y (n_59));
  NAND2X1 g12939(.A (\eps[14] [14]), .B (n_21), .Y (n_58));
  NAND2X1 g12940(.A (\eps[14] [10]), .B (n_48), .Y (n_57));
  OAI21X1 g3494(.A (\genblk1[15].inst_n_1114 ), .B (\eps[14] [13]), .C
       (\eps[14] [12]), .Y (n_56));
  NOR3X1 g12941(.A (1'b0), .B (1'b0), .C (n_39), .Y (n_55));
  NOR3X1 g12942(.A (1'b0), .B (1'b0), .C (n_40), .Y (n_51));
  OAI21X1 g12943(.A (query[2]), .B (query[3]), .C (n_4), .Y (n_50));
  OAI21X1 g12944(.A (n_24), .B (\eps[14] [14]), .C (n_21), .Y (n_54));
  OAI21X1 g12945(.A (n_32), .B (\eps[14] [6]), .C (n_22), .Y (n_53));
  AND2X1 g12946(.A (n_48), .B (n_44), .Y (n_52));
  OR2X1 g12947(.A (n_36), .B (result[15]), .Y (n_47));
  OR2X1 g12948(.A (\eps[14] [17]), .B (n_23), .Y (n_46));
  NAND2X1 g12949(.A (result[2]), .B (n_27), .Y (n_45));
  OR2X1 g12950(.A (\eps[14] [10]), .B (n_31), .Y (n_44));
  NAND2X1 g12951(.A (result[5]), .B (n_35), .Y (n_49));
  OR2X1 g12952(.A (\eps[14] [11]), .B (n_33), .Y (n_48));
  NAND2X1 g12953(.A (\genblk1[15].inst_n_1114 ), .B (\eps[14] [13]), .Y
       (n_42));
  NOR2X1 g12954(.A (1'b0), .B (1'b0), .Y (n_41));
  OR2X1 g12955(.A (1'b0), .B (1'b0), .Y (n_40));
  OR2X1 g12956(.A (1'b0), .B (1'b0), .Y (n_39));
  NOR2X1 g12957(.A (1'b0), .B (1'b0), .Y (n_38));
  NAND2X1 g12958(.A (result[13]), .B (n_34), .Y (n_43));
  NOR2X1 g12959(.A (\genblk1[15].inst_n_1114 ), .B (\eps[14] [13]), .Y
       (n_37));
  INVX1 g12960(.A (\eps[14] [17]), .Y (n_36));
  INVX1 g12961(.A (\eps[14] [7]), .Y (n_35));
  INVX1 g12962(.A (\eps[14] [15]), .Y (n_34));
  INVX1 g12963(.A (result[9]), .Y (n_33));
  INVX1 g12964(.A (result[4]), .Y (n_32));
  INVX1 g12965(.A (result[8]), .Y (n_31));
  INVX1 g12966(.A (result[6]), .Y (n_30));
  INVX1 g12967(.A (\eps[14] [8]), .Y (n_29));
  INVX1 g12968(.A (\eps[14] [5]), .Y (n_28));
  INVX1 g12969(.A (\eps[14] [4]), .Y (n_27));
  INVX1 g12970(.A (\eps[14] [9]), .Y (n_26));
  INVX1 g12971(.A (result[10]), .Y (n_25));
  INVX1 g12972(.A (result[12]), .Y (n_24));
  INVX1 g12973(.A (result[15]), .Y (n_23));
  BUFX2 drc_bufs3535(.A (n_74), .Y (n_20));
  BUFX2 drc_bufs3536(.A (n_79), .Y (n_19));
  BUFX2 drc_bufs3537(.A (n_41), .Y (n_18));
  BUFX2 drc_bufs3538(.A (n_37), .Y (n_17));
  BUFX2 drc_bufs3539(.A (n_78), .Y (n_16));
  BUFX2 drc_bufs3540(.A (n_38), .Y (n_15));
  BUFX2 drc_bufs3541(.A (n_42), .Y (n_14));
  BUFX2 drc_bufs3542(.A (n_57), .Y (n_13));
  BUFX2 drc_bufs3543(.A (n_58), .Y (n_12));
  BUFX2 drc_bufs3544(.A (n_87), .Y (n_11));
  BUFX2 drc_bufs3545(.A (n_67), .Y (n_10));
  BUFX2 drc_bufs3546(.A (n_65), .Y (n_9));
  BUFX2 drc_bufs3547(.A (n_59), .Y (n_8));
  BUFX2 drc_bufs3548(.A (n_88), .Y (n_7));
  BUFX2 drc_bufs12974(.A (n_77), .Y (n_6));
  BUFX2 drc_bufs3550(.A (n_76), .Y (n_5));
  BUFX2 drc_bufs12975(.A (n_45), .Y (n_4));
  BUFX2 drc_bufs12976(.A (n_84), .Y (n_3));
  BUFX2 drc_bufs12977(.A (n_80), .Y (n_2));
  BUFX2 drc_bufs12978(.A (n_85), .Y (n_1));
  BUFX2 drc_bufs12979(.A (n_90), .Y (\genblk1[15].inst_n_716 ));
  BUFX2 drc_bufs12980(.A (n_60), .Y (n_0));
  BUFX2 drc_bufs12981(.A (n_49), .Y (n_22));
  BUFX2 drc_bufs12982(.A (n_43), .Y (n_21));
  OR2X1 \genblk1[15].inst_SUB_UNS_OP_g1901 (.A (1'b0), .B (1'b0), .Y
       (\eps[15] [31]));
  INVX1 \genblk1[15].inst_SUB_UNS_OP_g1903 (.A
       (\genblk1[15].inst_SUB_UNS_OP_n_1034 ), .Y (\eps[15] [29]));
  NAND2X1 \genblk1[15].inst_SUB_UNS_OP_g1906 (.A
       (\genblk1[15].inst_SUB_UNS_OP_n_1030 ), .B (1'b1), .Y
       (\genblk1[15].inst_SUB_UNS_OP_n_893 ));
  NAND2X1 \genblk1[15].inst_SUB_UNS_OP_g1908 (.A (1'b0), .B (1'b1), .Y
       (\genblk1[15].inst_SUB_UNS_OP_n_898 ));
  INVX1 \genblk1[15].inst_SUB_UNS_OP_g1912 (.A
       (\genblk1[15].inst_SUB_UNS_OP_n_1033 ), .Y (\eps[15] [26]));
  NAND2X1 \genblk1[15].inst_SUB_UNS_OP_g1915 (.A
       (\genblk1[15].inst_SUB_UNS_OP_n_1026 ), .B (1'b1), .Y
       (\genblk1[15].inst_SUB_UNS_OP_n_909 ));
  NAND2X1 \genblk1[15].inst_SUB_UNS_OP_g1916 (.A (1'b0), .B (1'b1), .Y
       (\genblk1[15].inst_SUB_UNS_OP_n_911 ));
  INVX1 \genblk1[15].inst_SUB_UNS_OP_g1921 (.A
       (\genblk1[15].inst_SUB_UNS_OP_n_1031 ), .Y (\eps[15] [23]));
  INVX1 \genblk1[15].inst_SUB_UNS_OP_g1930 (.A
       (\genblk1[15].inst_SUB_UNS_OP_n_1032 ), .Y (\eps[15] [20]));
  NAND2X1 \genblk1[15].inst_SUB_UNS_OP_g1933 (.A
       (\genblk1[15].inst_SUB_UNS_OP_n_1028 ), .B (1'b1), .Y
       (\genblk1[15].inst_SUB_UNS_OP_n_941 ));
  NAND2X1 \genblk1[15].inst_SUB_UNS_OP_g1934 (.A (1'b0), .B (1'b1), .Y
       (\genblk1[15].inst_SUB_UNS_OP_n_943 ));
  NAND2X1 \genblk1[15].inst_SUB_UNS_OP_g1936 (.A
       (\genblk1[15].inst_SUB_UNS_OP_n_1029 ), .B (1'b1), .Y
       (\genblk1[15].inst_SUB_UNS_OP_n_948 ));
  NAND2X1 \genblk1[15].inst_SUB_UNS_OP_g1937 (.A (\eps[14] [18]), .B
       (\genblk1[15].inst_SUB_UNS_OP_n_954 ), .Y
       (\genblk1[15].inst_SUB_UNS_OP_n_949 ));
  FAX1 \genblk1[15].inst_SUB_UNS_OP_g1939 (.A (\eps[14] [17]), .B
       (\genblk1[15].inst_SUB_UNS_OP_n_994 ), .C
       (\genblk1[15].inst_SUB_UNS_OP_n_957 ), .YC
       (\genblk1[15].inst_SUB_UNS_OP_n_954 ), .YS (\eps[15] [17]));
  FAX1 \genblk1[15].inst_SUB_UNS_OP_g1940 (.A (\eps[14] [16]), .B
       (\genblk1[15].inst_SUB_UNS_OP_n_1017 ), .C
       (\genblk1[15].inst_SUB_UNS_OP_n_959 ), .YC
       (\genblk1[15].inst_SUB_UNS_OP_n_957 ), .YS (\eps[15] [16]));
  FAX1 \genblk1[15].inst_SUB_UNS_OP_g1941 (.A (\eps[14] [15]), .B
       (\genblk1[15].inst_SUB_UNS_OP_n_1012 ), .C
       (\genblk1[15].inst_SUB_UNS_OP_n_961 ), .YC
       (\genblk1[15].inst_SUB_UNS_OP_n_959 ), .YS (\eps[15] [15]));
  FAX1 \genblk1[15].inst_SUB_UNS_OP_g1942 (.A (\eps[14] [14]), .B
       (\genblk1[15].inst_SUB_UNS_OP_n_1008 ), .C
       (\genblk1[15].inst_SUB_UNS_OP_n_963 ), .YC
       (\genblk1[15].inst_SUB_UNS_OP_n_961 ), .YS (\eps[15] [14]));
  FAX1 \genblk1[15].inst_SUB_UNS_OP_g1943 (.A (\eps[14] [13]), .B
       (\genblk1[15].inst_SUB_UNS_OP_n_1018 ), .C
       (\genblk1[15].inst_SUB_UNS_OP_n_965 ), .YC
       (\genblk1[15].inst_SUB_UNS_OP_n_963 ), .YS (\eps[15] [13]));
  FAX1 \genblk1[15].inst_SUB_UNS_OP_g1944 (.A (\eps[14] [12]), .B
       (\genblk1[15].inst_SUB_UNS_OP_n_991 ), .C
       (\genblk1[15].inst_SUB_UNS_OP_n_967 ), .YC
       (\genblk1[15].inst_SUB_UNS_OP_n_965 ), .YS (\eps[15] [12]));
  FAX1 \genblk1[15].inst_SUB_UNS_OP_g1945 (.A (\eps[14] [11]), .B
       (\genblk1[15].inst_SUB_UNS_OP_n_1007 ), .C
       (\genblk1[15].inst_SUB_UNS_OP_n_969 ), .YC
       (\genblk1[15].inst_SUB_UNS_OP_n_967 ), .YS (\eps[15] [11]));
  FAX1 \genblk1[15].inst_SUB_UNS_OP_g1946 (.A (\eps[14] [10]), .B
       (\genblk1[15].inst_SUB_UNS_OP_n_1016 ), .C
       (\genblk1[15].inst_SUB_UNS_OP_n_971 ), .YC
       (\genblk1[15].inst_SUB_UNS_OP_n_969 ), .YS (\eps[15] [10]));
  FAX1 \genblk1[15].inst_SUB_UNS_OP_g1947 (.A (\eps[14] [9]), .B
       (\genblk1[15].inst_SUB_UNS_OP_n_993 ), .C
       (\genblk1[15].inst_SUB_UNS_OP_n_973 ), .YC
       (\genblk1[15].inst_SUB_UNS_OP_n_971 ), .YS (\eps[15] [9]));
  FAX1 \genblk1[15].inst_SUB_UNS_OP_g1948 (.A (\eps[14] [8]), .B
       (\genblk1[15].inst_SUB_UNS_OP_n_1019 ), .C
       (\genblk1[15].inst_SUB_UNS_OP_n_975 ), .YC
       (\genblk1[15].inst_SUB_UNS_OP_n_973 ), .YS (\eps[15] [8]));
  FAX1 \genblk1[15].inst_SUB_UNS_OP_g1949 (.A (\eps[14] [7]), .B
       (\genblk1[15].inst_SUB_UNS_OP_n_999 ), .C
       (\genblk1[15].inst_SUB_UNS_OP_n_977 ), .YC
       (\genblk1[15].inst_SUB_UNS_OP_n_975 ), .YS (\eps[15] [7]));
  FAX1 \genblk1[15].inst_SUB_UNS_OP_g1950 (.A (\eps[14] [6]), .B
       (\genblk1[15].inst_SUB_UNS_OP_n_1004 ), .C
       (\genblk1[15].inst_SUB_UNS_OP_n_979 ), .YC
       (\genblk1[15].inst_SUB_UNS_OP_n_977 ), .YS (\eps[15] [6]));
  FAX1 \genblk1[15].inst_SUB_UNS_OP_g1951 (.A (\eps[14] [5]), .B
       (\genblk1[15].inst_SUB_UNS_OP_n_1011 ), .C
       (\genblk1[15].inst_SUB_UNS_OP_n_981 ), .YC
       (\genblk1[15].inst_SUB_UNS_OP_n_979 ), .YS (\eps[15] [5]));
  FAX1 \genblk1[15].inst_SUB_UNS_OP_g1952 (.A (\eps[14] [4]), .B
       (\genblk1[15].inst_SUB_UNS_OP_n_990 ), .C
       (\genblk1[15].inst_SUB_UNS_OP_n_983 ), .YC
       (\genblk1[15].inst_SUB_UNS_OP_n_981 ), .YS (\eps[15] [4]));
  INVX1 \genblk1[15].inst_SUB_UNS_OP_g1953 (.A
       (\genblk1[15].inst_SUB_UNS_OP_n_984 ), .Y (\eps[15] [3]));
  INVX1 \genblk1[15].inst_SUB_UNS_OP_g1954 (.A
       (\genblk1[15].inst_SUB_UNS_OP_n_985 ), .Y
       (\genblk1[15].inst_SUB_UNS_OP_n_983 ));
  HAX1 \genblk1[15].inst_SUB_UNS_OP_g1955 (.A
       (\genblk1[15].inst_SUB_UNS_OP_n_998 ), .B
       (\genblk1[15].inst_SUB_UNS_OP_n_988 ), .YC
       (\genblk1[15].inst_SUB_UNS_OP_n_985 ), .YS
       (\genblk1[15].inst_SUB_UNS_OP_n_984 ));
  INVX1 \genblk1[15].inst_SUB_UNS_OP_g1956 (.A
       (\genblk1[15].inst_SUB_UNS_OP_n_987 ), .Y (\eps[15] [2]));
  HAX1 \genblk1[15].inst_SUB_UNS_OP_g1957 (.A
       (\genblk1[15].inst_SUB_UNS_OP_n_992 ), .B (result[1]), .YC
       (\genblk1[15].inst_SUB_UNS_OP_n_988 ), .YS
       (\genblk1[15].inst_SUB_UNS_OP_n_987 ));
  INVX1 \genblk1[15].inst_SUB_UNS_OP_g1958 (.A (\genblk1[15].inst_n_725
       ), .Y (\genblk1[15].inst_SUB_UNS_OP_n_990 ));
  INVX1 \genblk1[15].inst_SUB_UNS_OP_g1959 (.A (\genblk1[15].inst_n_717
       ), .Y (\genblk1[15].inst_SUB_UNS_OP_n_991 ));
  INVX1 \genblk1[15].inst_SUB_UNS_OP_g1960 (.A (query[2]), .Y
       (\genblk1[15].inst_SUB_UNS_OP_n_992 ));
  INVX1 \genblk1[15].inst_SUB_UNS_OP_g1961 (.A (\genblk1[15].inst_n_720
       ), .Y (\genblk1[15].inst_SUB_UNS_OP_n_993 ));
  INVX1 \genblk1[15].inst_SUB_UNS_OP_g1962 (.A (\genblk1[15].inst_n_712
       ), .Y (\genblk1[15].inst_SUB_UNS_OP_n_994 ));
  INVX1 \genblk1[15].inst_SUB_UNS_OP_g1963 (.A (query[3]), .Y
       (\genblk1[15].inst_SUB_UNS_OP_n_998 ));
  INVX1 \genblk1[15].inst_SUB_UNS_OP_g1964 (.A (\genblk1[15].inst_n_722
       ), .Y (\genblk1[15].inst_SUB_UNS_OP_n_999 ));
  INVX1 \genblk1[15].inst_SUB_UNS_OP_g1965 (.A (\genblk1[15].inst_n_723
       ), .Y (\genblk1[15].inst_SUB_UNS_OP_n_1004 ));
  INVX1 \genblk1[15].inst_SUB_UNS_OP_g1967 (.A (\genblk1[15].inst_n_718
       ), .Y (\genblk1[15].inst_SUB_UNS_OP_n_1007 ));
  INVX1 \genblk1[15].inst_SUB_UNS_OP_g1968 (.A (\genblk1[15].inst_n_715
       ), .Y (\genblk1[15].inst_SUB_UNS_OP_n_1008 ));
  INVX1 \genblk1[15].inst_SUB_UNS_OP_g1970 (.A (\genblk1[15].inst_n_724
       ), .Y (\genblk1[15].inst_SUB_UNS_OP_n_1011 ));
  INVX1 \genblk1[15].inst_SUB_UNS_OP_g1971 (.A (\genblk1[15].inst_n_714
       ), .Y (\genblk1[15].inst_SUB_UNS_OP_n_1012 ));
  INVX1 \genblk1[15].inst_SUB_UNS_OP_g1973 (.A (\genblk1[15].inst_n_719
       ), .Y (\genblk1[15].inst_SUB_UNS_OP_n_1016 ));
  INVX1 \genblk1[15].inst_SUB_UNS_OP_g1974 (.A (\genblk1[15].inst_n_713
       ), .Y (\genblk1[15].inst_SUB_UNS_OP_n_1017 ));
  INVX1 \genblk1[15].inst_SUB_UNS_OP_g1975 (.A (\genblk1[15].inst_n_716
       ), .Y (\genblk1[15].inst_SUB_UNS_OP_n_1018 ));
  INVX1 \genblk1[15].inst_SUB_UNS_OP_g1976 (.A (\genblk1[15].inst_n_721
       ), .Y (\genblk1[15].inst_SUB_UNS_OP_n_1019 ));
  BUFX2 \genblk1[15].inst_SUB_UNS_OP_drc_bufs (.A
       (\genblk1[15].inst_SUB_UNS_OP_n_893 ), .Y (\eps[15] [28]));
  BUFX2 \genblk1[15].inst_SUB_UNS_OP_drc_bufs1977 (.A
       (\genblk1[15].inst_SUB_UNS_OP_n_909 ), .Y (\eps[15] [25]));
  BUFX2 \genblk1[15].inst_SUB_UNS_OP_drc_bufs1978 (.A
       (\genblk1[15].inst_SUB_UNS_OP_n_941 ), .Y (\eps[15] [19]));
  BUFX2 \genblk1[15].inst_SUB_UNS_OP_drc_bufs1979 (.A
       (\genblk1[15].inst_SUB_UNS_OP_n_948 ), .Y (\eps[15] [18]));
  BUFX2 \genblk1[15].inst_SUB_UNS_OP_drc_bufs1981 (.A
       (\genblk1[15].inst_SUB_UNS_OP_n_911 ), .Y
       (\genblk1[15].inst_SUB_UNS_OP_n_1026 ));
  BUFX2 \genblk1[15].inst_SUB_UNS_OP_drc_bufs1983 (.A
       (\genblk1[15].inst_SUB_UNS_OP_n_943 ), .Y
       (\genblk1[15].inst_SUB_UNS_OP_n_1028 ));
  BUFX2 \genblk1[15].inst_SUB_UNS_OP_drc_bufs1984 (.A
       (\genblk1[15].inst_SUB_UNS_OP_n_949 ), .Y
       (\genblk1[15].inst_SUB_UNS_OP_n_1029 ));
  BUFX2 \genblk1[15].inst_SUB_UNS_OP_drc_bufs1985 (.A
       (\genblk1[15].inst_SUB_UNS_OP_n_898 ), .Y
       (\genblk1[15].inst_SUB_UNS_OP_n_1030 ));
  BUFX2 \genblk1[15].inst_SUB_UNS_OP_drc_bufs1986 (.A (1'b1), .Y
       (\genblk1[15].inst_SUB_UNS_OP_n_1031 ));
  BUFX2 \genblk1[15].inst_SUB_UNS_OP_drc_bufs1987 (.A (1'b1), .Y
       (\genblk1[15].inst_SUB_UNS_OP_n_1032 ));
  BUFX2 \genblk1[15].inst_SUB_UNS_OP_drc_bufs1988 (.A (1'b1), .Y
       (\genblk1[15].inst_SUB_UNS_OP_n_1033 ));
  BUFX2 \genblk1[15].inst_SUB_UNS_OP_drc_bufs1989 (.A (1'b1), .Y
       (\genblk1[15].inst_SUB_UNS_OP_n_1034 ));
  XNOR2X1 \genblk1[14].inst_SUB_UNS_OP_g1801 (.A
       (\genblk1[14].inst_SUB_UNS_OP_n_909 ), .B
       (\genblk1[14].inst_SUB_UNS_OP_n_940 ), .Y (\eps[14] [18]));
  FAX1 \genblk1[14].inst_SUB_UNS_OP_g1803 (.A (\eps[13] [17]), .B
       (\genblk1[14].inst_SUB_UNS_OP_n_949 ), .C
       (\genblk1[14].inst_SUB_UNS_OP_n_912 ), .YC
       (\genblk1[14].inst_SUB_UNS_OP_n_909 ), .YS (\eps[14] [17]));
  FAX1 \genblk1[14].inst_SUB_UNS_OP_g1804 (.A (\eps[13] [16]), .B
       (\genblk1[14].inst_SUB_UNS_OP_n_955 ), .C
       (\genblk1[14].inst_SUB_UNS_OP_n_914 ), .YC
       (\genblk1[14].inst_SUB_UNS_OP_n_912 ), .YS (\eps[14] [16]));
  FAX1 \genblk1[14].inst_SUB_UNS_OP_g1805 (.A (\eps[13] [15]), .B
       (\genblk1[14].inst_SUB_UNS_OP_n_961 ), .C
       (\genblk1[14].inst_SUB_UNS_OP_n_916 ), .YC
       (\genblk1[14].inst_SUB_UNS_OP_n_914 ), .YS (\eps[14] [15]));
  FAX1 \genblk1[14].inst_SUB_UNS_OP_g1806 (.A (\eps[13] [14]), .B
       (\genblk1[14].inst_SUB_UNS_OP_n_951 ), .C
       (\genblk1[14].inst_SUB_UNS_OP_n_918 ), .YC
       (\genblk1[14].inst_SUB_UNS_OP_n_916 ), .YS (\eps[14] [14]));
  FAX1 \genblk1[14].inst_SUB_UNS_OP_g1807 (.A (\eps[13] [13]), .B
       (\genblk1[14].inst_SUB_UNS_OP_n_945 ), .C
       (\genblk1[14].inst_SUB_UNS_OP_n_920 ), .YC
       (\genblk1[14].inst_SUB_UNS_OP_n_918 ), .YS (\eps[14] [13]));
  FAX1 \genblk1[14].inst_SUB_UNS_OP_g1808 (.A (\eps[13] [12]), .B
       (\genblk1[14].inst_SUB_UNS_OP_n_968 ), .C
       (\genblk1[14].inst_SUB_UNS_OP_n_922 ), .YC
       (\genblk1[14].inst_SUB_UNS_OP_n_920 ), .YS (\eps[14] [12]));
  FAX1 \genblk1[14].inst_SUB_UNS_OP_g1809 (.A (\eps[13] [11]), .B
       (\genblk1[14].inst_SUB_UNS_OP_n_966 ), .C
       (\genblk1[14].inst_SUB_UNS_OP_n_924 ), .YC
       (\genblk1[14].inst_SUB_UNS_OP_n_922 ), .YS (\eps[14] [11]));
  FAX1 \genblk1[14].inst_SUB_UNS_OP_g1810 (.A (\eps[13] [10]), .B
       (\genblk1[14].inst_SUB_UNS_OP_n_959 ), .C
       (\genblk1[14].inst_SUB_UNS_OP_n_926 ), .YC
       (\genblk1[14].inst_SUB_UNS_OP_n_924 ), .YS (\eps[14] [10]));
  FAX1 \genblk1[14].inst_SUB_UNS_OP_g1811 (.A (\eps[13] [9]), .B
       (\genblk1[14].inst_SUB_UNS_OP_n_950 ), .C
       (\genblk1[14].inst_SUB_UNS_OP_n_928 ), .YC
       (\genblk1[14].inst_SUB_UNS_OP_n_926 ), .YS (\eps[14] [9]));
  FAX1 \genblk1[14].inst_SUB_UNS_OP_g1812 (.A (\eps[13] [8]), .B
       (\genblk1[14].inst_SUB_UNS_OP_n_972 ), .C
       (\genblk1[14].inst_SUB_UNS_OP_n_930 ), .YC
       (\genblk1[14].inst_SUB_UNS_OP_n_928 ), .YS (\eps[14] [8]));
  FAX1 \genblk1[14].inst_SUB_UNS_OP_g1813 (.A (\eps[13] [7]), .B
       (\genblk1[14].inst_SUB_UNS_OP_n_947 ), .C
       (\genblk1[14].inst_SUB_UNS_OP_n_932 ), .YC
       (\genblk1[14].inst_SUB_UNS_OP_n_930 ), .YS (\eps[14] [7]));
  FAX1 \genblk1[14].inst_SUB_UNS_OP_g1814 (.A (\eps[13] [6]), .B
       (\genblk1[14].inst_SUB_UNS_OP_n_952 ), .C
       (\genblk1[14].inst_SUB_UNS_OP_n_934 ), .YC
       (\genblk1[14].inst_SUB_UNS_OP_n_932 ), .YS (\eps[14] [6]));
  INVX1 \genblk1[14].inst_SUB_UNS_OP_g1815 (.A
       (\genblk1[14].inst_SUB_UNS_OP_n_935 ), .Y (\eps[14] [5]));
  INVX1 \genblk1[14].inst_SUB_UNS_OP_g1816 (.A
       (\genblk1[14].inst_SUB_UNS_OP_n_936 ), .Y
       (\genblk1[14].inst_SUB_UNS_OP_n_934 ));
  HAX1 \genblk1[14].inst_SUB_UNS_OP_g1817 (.A
       (\genblk1[14].inst_SUB_UNS_OP_n_956 ), .B
       (\genblk1[14].inst_SUB_UNS_OP_n_939 ), .YC
       (\genblk1[14].inst_SUB_UNS_OP_n_936 ), .YS
       (\genblk1[14].inst_SUB_UNS_OP_n_935 ));
  INVX1 \genblk1[14].inst_SUB_UNS_OP_g1818 (.A
       (\genblk1[14].inst_SUB_UNS_OP_n_938 ), .Y (\eps[14] [4]));
  HAX1 \genblk1[14].inst_SUB_UNS_OP_g1819 (.A
       (\genblk1[14].inst_SUB_UNS_OP_n_960 ), .B (result[2]), .YC
       (\genblk1[14].inst_SUB_UNS_OP_n_939 ), .YS
       (\genblk1[14].inst_SUB_UNS_OP_n_938 ));
  OR2X1 \genblk1[14].inst_SUB_UNS_OP_g1820 (.A
       (\genblk1[14].inst_SUB_UNS_OP_n_941 ), .B
       (\genblk1[14].inst_SUB_UNS_OP_n_943 ), .Y
       (\genblk1[14].inst_SUB_UNS_OP_n_940 ));
  AND2X1 \genblk1[14].inst_SUB_UNS_OP_g1821 (.A
       (\genblk1[14].inst_SUB_UNS_OP_n_953 ), .B (\eps[13] [18]), .Y
       (\genblk1[14].inst_SUB_UNS_OP_n_941 ));
  AND2X1 \genblk1[14].inst_SUB_UNS_OP_g1823 (.A
       (\genblk1[14].inst_n_711 ), .B
       (\genblk1[14].inst_SUB_UNS_OP_n_964 ), .Y
       (\genblk1[14].inst_SUB_UNS_OP_n_943 ));
  INVX1 \genblk1[14].inst_SUB_UNS_OP_g1825 (.A (\genblk1[14].inst_n_716
       ), .Y (\genblk1[14].inst_SUB_UNS_OP_n_945 ));
  INVX1 \genblk1[14].inst_SUB_UNS_OP_g1827 (.A (\genblk1[14].inst_n_722
       ), .Y (\genblk1[14].inst_SUB_UNS_OP_n_947 ));
  INVX1 \genblk1[14].inst_SUB_UNS_OP_g1829 (.A (\genblk1[14].inst_n_712
       ), .Y (\genblk1[14].inst_SUB_UNS_OP_n_949 ));
  INVX1 \genblk1[14].inst_SUB_UNS_OP_g1830 (.A (\genblk1[14].inst_n_720
       ), .Y (\genblk1[14].inst_SUB_UNS_OP_n_950 ));
  INVX1 \genblk1[14].inst_SUB_UNS_OP_g1831 (.A (\genblk1[14].inst_n_715
       ), .Y (\genblk1[14].inst_SUB_UNS_OP_n_951 ));
  INVX1 \genblk1[14].inst_SUB_UNS_OP_g1832 (.A (\genblk1[14].inst_n_723
       ), .Y (\genblk1[14].inst_SUB_UNS_OP_n_952 ));
  INVX1 \genblk1[14].inst_SUB_UNS_OP_g1833 (.A (\genblk1[14].inst_n_711
       ), .Y (\genblk1[14].inst_SUB_UNS_OP_n_953 ));
  INVX1 \genblk1[14].inst_SUB_UNS_OP_g1834 (.A (\genblk1[14].inst_n_713
       ), .Y (\genblk1[14].inst_SUB_UNS_OP_n_955 ));
  INVX1 \genblk1[14].inst_SUB_UNS_OP_g1835 (.A (query[5]), .Y
       (\genblk1[14].inst_SUB_UNS_OP_n_956 ));
  INVX1 \genblk1[14].inst_SUB_UNS_OP_g1837 (.A (\genblk1[14].inst_n_719
       ), .Y (\genblk1[14].inst_SUB_UNS_OP_n_959 ));
  INVX1 \genblk1[14].inst_SUB_UNS_OP_g1838 (.A (query[4]), .Y
       (\genblk1[14].inst_SUB_UNS_OP_n_960 ));
  INVX1 \genblk1[14].inst_SUB_UNS_OP_g1839 (.A (\genblk1[14].inst_n_714
       ), .Y (\genblk1[14].inst_SUB_UNS_OP_n_961 ));
  INVX1 \genblk1[14].inst_SUB_UNS_OP_g1842 (.A (\eps[13] [18]), .Y
       (\genblk1[14].inst_SUB_UNS_OP_n_964 ));
  INVX1 \genblk1[14].inst_SUB_UNS_OP_g1843 (.A (\genblk1[14].inst_n_718
       ), .Y (\genblk1[14].inst_SUB_UNS_OP_n_966 ));
  INVX1 \genblk1[14].inst_SUB_UNS_OP_g1844 (.A (\genblk1[14].inst_n_717
       ), .Y (\genblk1[14].inst_SUB_UNS_OP_n_968 ));
  INVX1 \genblk1[14].inst_SUB_UNS_OP_g1848 (.A (\genblk1[14].inst_n_721
       ), .Y (\genblk1[14].inst_SUB_UNS_OP_n_972 ));
  INVX1 \genblk1[13].inst_SUB_UNS_OP_g1660 (.A
       (\genblk1[13].inst_SUB_UNS_OP_n_927 ), .Y (\eps[13] [24]));
  FAX1 \genblk1[13].inst_SUB_UNS_OP_g1674 (.A (\eps[12] [19]), .B
       (\genblk1[13].inst_SUB_UNS_OP_n_901 ), .C
       (\genblk1[13].inst_SUB_UNS_OP_n_872 ), .YC
       (\genblk1[13].inst_SUB_UNS_OP_n_869 ), .YS (\eps[13] [19]));
  FAX1 \genblk1[13].inst_SUB_UNS_OP_g1675 (.A (\eps[12] [18]), .B
       (\genblk1[13].inst_SUB_UNS_OP_n_919 ), .C
       (\genblk1[13].inst_SUB_UNS_OP_n_874 ), .YC
       (\genblk1[13].inst_SUB_UNS_OP_n_872 ), .YS (\eps[13] [18]));
  FAX1 \genblk1[13].inst_SUB_UNS_OP_g1676 (.A (\eps[12] [17]), .B
       (\genblk1[13].inst_SUB_UNS_OP_n_907 ), .C
       (\genblk1[13].inst_SUB_UNS_OP_n_876 ), .YC
       (\genblk1[13].inst_SUB_UNS_OP_n_874 ), .YS (\eps[13] [17]));
  FAX1 \genblk1[13].inst_SUB_UNS_OP_g1677 (.A (\eps[12] [16]), .B
       (\genblk1[13].inst_SUB_UNS_OP_n_902 ), .C
       (\genblk1[13].inst_SUB_UNS_OP_n_878 ), .YC
       (\genblk1[13].inst_SUB_UNS_OP_n_876 ), .YS (\eps[13] [16]));
  FAX1 \genblk1[13].inst_SUB_UNS_OP_g1678 (.A (\eps[12] [15]), .B
       (\genblk1[13].inst_SUB_UNS_OP_n_905 ), .C
       (\genblk1[13].inst_SUB_UNS_OP_n_880 ), .YC
       (\genblk1[13].inst_SUB_UNS_OP_n_878 ), .YS (\eps[13] [15]));
  FAX1 \genblk1[13].inst_SUB_UNS_OP_g1679 (.A (\eps[12] [14]), .B
       (\genblk1[13].inst_SUB_UNS_OP_n_906 ), .C
       (\genblk1[13].inst_SUB_UNS_OP_n_882 ), .YC
       (\genblk1[13].inst_SUB_UNS_OP_n_880 ), .YS (\eps[13] [14]));
  FAX1 \genblk1[13].inst_SUB_UNS_OP_g1680 (.A (\eps[12] [13]), .B
       (\genblk1[13].inst_SUB_UNS_OP_n_904 ), .C
       (\genblk1[13].inst_SUB_UNS_OP_n_884 ), .YC
       (\genblk1[13].inst_SUB_UNS_OP_n_882 ), .YS (\eps[13] [13]));
  FAX1 \genblk1[13].inst_SUB_UNS_OP_g1681 (.A (\eps[12] [12]), .B
       (\genblk1[13].inst_SUB_UNS_OP_n_911 ), .C
       (\genblk1[13].inst_SUB_UNS_OP_n_886 ), .YC
       (\genblk1[13].inst_SUB_UNS_OP_n_884 ), .YS (\eps[13] [12]));
  FAX1 \genblk1[13].inst_SUB_UNS_OP_g1682 (.A (\eps[12] [11]), .B
       (\genblk1[13].inst_SUB_UNS_OP_n_920 ), .C
       (\genblk1[13].inst_SUB_UNS_OP_n_888 ), .YC
       (\genblk1[13].inst_SUB_UNS_OP_n_886 ), .YS (\eps[13] [11]));
  FAX1 \genblk1[13].inst_SUB_UNS_OP_g1683 (.A (\eps[12] [10]), .B
       (\genblk1[13].inst_SUB_UNS_OP_n_921 ), .C
       (\genblk1[13].inst_SUB_UNS_OP_n_890 ), .YC
       (\genblk1[13].inst_SUB_UNS_OP_n_888 ), .YS (\eps[13] [10]));
  FAX1 \genblk1[13].inst_SUB_UNS_OP_g1684 (.A (\eps[12] [9]), .B
       (\genblk1[13].inst_SUB_UNS_OP_n_916 ), .C
       (\genblk1[13].inst_SUB_UNS_OP_n_892 ), .YC
       (\genblk1[13].inst_SUB_UNS_OP_n_890 ), .YS (\eps[13] [9]));
  FAX1 \genblk1[13].inst_SUB_UNS_OP_g1685 (.A (\eps[12] [8]), .B
       (\genblk1[13].inst_SUB_UNS_OP_n_923 ), .C
       (\genblk1[13].inst_SUB_UNS_OP_n_894 ), .YC
       (\genblk1[13].inst_SUB_UNS_OP_n_892 ), .YS (\eps[13] [8]));
  INVX1 \genblk1[13].inst_SUB_UNS_OP_g1686 (.A
       (\genblk1[13].inst_SUB_UNS_OP_n_895 ), .Y (\eps[13] [7]));
  INVX1 \genblk1[13].inst_SUB_UNS_OP_g1687 (.A
       (\genblk1[13].inst_SUB_UNS_OP_n_896 ), .Y
       (\genblk1[13].inst_SUB_UNS_OP_n_894 ));
  HAX1 \genblk1[13].inst_SUB_UNS_OP_g1688 (.A
       (\genblk1[13].inst_SUB_UNS_OP_n_924 ), .B
       (\genblk1[13].inst_SUB_UNS_OP_n_899 ), .YC
       (\genblk1[13].inst_SUB_UNS_OP_n_896 ), .YS
       (\genblk1[13].inst_SUB_UNS_OP_n_895 ));
  INVX1 \genblk1[13].inst_SUB_UNS_OP_g1689 (.A
       (\genblk1[13].inst_SUB_UNS_OP_n_898 ), .Y (\eps[13] [6]));
  HAX1 \genblk1[13].inst_SUB_UNS_OP_g1690 (.A
       (\genblk1[13].inst_SUB_UNS_OP_n_903 ), .B (result[3]), .YC
       (\genblk1[13].inst_SUB_UNS_OP_n_899 ), .YS
       (\genblk1[13].inst_SUB_UNS_OP_n_898 ));
  INVX1 \genblk1[13].inst_SUB_UNS_OP_g1691 (.A (\genblk1[13].inst_n_710
       ), .Y (\genblk1[13].inst_SUB_UNS_OP_n_901 ));
  INVX1 \genblk1[13].inst_SUB_UNS_OP_g1692 (.A (\genblk1[13].inst_n_713
       ), .Y (\genblk1[13].inst_SUB_UNS_OP_n_902 ));
  INVX1 \genblk1[13].inst_SUB_UNS_OP_g1693 (.A (query[6]), .Y
       (\genblk1[13].inst_SUB_UNS_OP_n_903 ));
  INVX1 \genblk1[13].inst_SUB_UNS_OP_g1694 (.A (\genblk1[13].inst_n_716
       ), .Y (\genblk1[13].inst_SUB_UNS_OP_n_904 ));
  INVX1 \genblk1[13].inst_SUB_UNS_OP_g1695 (.A (\genblk1[13].inst_n_714
       ), .Y (\genblk1[13].inst_SUB_UNS_OP_n_905 ));
  INVX1 \genblk1[13].inst_SUB_UNS_OP_g1696 (.A (\genblk1[13].inst_n_715
       ), .Y (\genblk1[13].inst_SUB_UNS_OP_n_906 ));
  INVX1 \genblk1[13].inst_SUB_UNS_OP_g1697 (.A (\genblk1[13].inst_n_712
       ), .Y (\genblk1[13].inst_SUB_UNS_OP_n_907 ));
  INVX1 \genblk1[13].inst_SUB_UNS_OP_g1699 (.A (\genblk1[13].inst_n_717
       ), .Y (\genblk1[13].inst_SUB_UNS_OP_n_911 ));
  INVX1 \genblk1[13].inst_SUB_UNS_OP_g1700 (.A (\genblk1[13].inst_n_720
       ), .Y (\genblk1[13].inst_SUB_UNS_OP_n_916 ));
  INVX1 \genblk1[13].inst_SUB_UNS_OP_g1702 (.A (\genblk1[13].inst_n_711
       ), .Y (\genblk1[13].inst_SUB_UNS_OP_n_919 ));
  INVX1 \genblk1[13].inst_SUB_UNS_OP_g1703 (.A (\genblk1[13].inst_n_718
       ), .Y (\genblk1[13].inst_SUB_UNS_OP_n_920 ));
  INVX1 \genblk1[13].inst_SUB_UNS_OP_g1704 (.A (\genblk1[13].inst_n_719
       ), .Y (\genblk1[13].inst_SUB_UNS_OP_n_921 ));
  INVX1 \genblk1[13].inst_SUB_UNS_OP_g1705 (.A (\genblk1[13].inst_n_721
       ), .Y (\genblk1[13].inst_SUB_UNS_OP_n_923 ));
  INVX1 \genblk1[13].inst_SUB_UNS_OP_g1706 (.A (query[7]), .Y
       (\genblk1[13].inst_SUB_UNS_OP_n_924 ));
  BUFX2 \genblk1[13].inst_SUB_UNS_OP_drc_bufs1708 (.A (1'b1), .Y
       (\genblk1[13].inst_SUB_UNS_OP_n_927 ));
  OR2X1 \genblk1[12].inst_SUB_UNS_OP_g1531 (.A (1'b0), .B (1'b0), .Y
       (\eps[12] [31]));
  XNOR2X1 \genblk1[12].inst_SUB_UNS_OP_g1550 (.A
       (\genblk1[12].inst_SUB_UNS_OP_n_822 ), .B
       (\genblk1[12].inst_SUB_UNS_OP_n_849 ), .Y (\eps[12] [20]));
  FAX1 \genblk1[12].inst_SUB_UNS_OP_g1552 (.A (\eps[11] [19]), .B
       (\genblk1[12].inst_SUB_UNS_OP_n_853 ), .C
       (\genblk1[12].inst_SUB_UNS_OP_n_825 ), .YC
       (\genblk1[12].inst_SUB_UNS_OP_n_822 ), .YS (\eps[12] [19]));
  FAX1 \genblk1[12].inst_SUB_UNS_OP_g1553 (.A (\eps[11] [18]), .B
       (\genblk1[12].inst_SUB_UNS_OP_n_859 ), .C
       (\genblk1[12].inst_SUB_UNS_OP_n_827 ), .YC
       (\genblk1[12].inst_SUB_UNS_OP_n_825 ), .YS (\eps[12] [18]));
  FAX1 \genblk1[12].inst_SUB_UNS_OP_g1554 (.A (\eps[11] [17]), .B
       (\genblk1[12].inst_SUB_UNS_OP_n_862 ), .C
       (\genblk1[12].inst_SUB_UNS_OP_n_829 ), .YC
       (\genblk1[12].inst_SUB_UNS_OP_n_827 ), .YS (\eps[12] [17]));
  FAX1 \genblk1[12].inst_SUB_UNS_OP_g1555 (.A (\eps[11] [16]), .B
       (\genblk1[12].inst_SUB_UNS_OP_n_857 ), .C
       (\genblk1[12].inst_SUB_UNS_OP_n_831 ), .YC
       (\genblk1[12].inst_SUB_UNS_OP_n_829 ), .YS (\eps[12] [16]));
  FAX1 \genblk1[12].inst_SUB_UNS_OP_g1556 (.A (\eps[11] [15]), .B
       (\genblk1[12].inst_SUB_UNS_OP_n_866 ), .C
       (\genblk1[12].inst_SUB_UNS_OP_n_833 ), .YC
       (\genblk1[12].inst_SUB_UNS_OP_n_831 ), .YS (\eps[12] [15]));
  FAX1 \genblk1[12].inst_SUB_UNS_OP_g1557 (.A (\eps[11] [14]), .B
       (\genblk1[12].inst_SUB_UNS_OP_n_874 ), .C
       (\genblk1[12].inst_SUB_UNS_OP_n_835 ), .YC
       (\genblk1[12].inst_SUB_UNS_OP_n_833 ), .YS (\eps[12] [14]));
  FAX1 \genblk1[12].inst_SUB_UNS_OP_g1558 (.A (\eps[11] [13]), .B
       (\genblk1[12].inst_SUB_UNS_OP_n_873 ), .C
       (\genblk1[12].inst_SUB_UNS_OP_n_837 ), .YC
       (\genblk1[12].inst_SUB_UNS_OP_n_835 ), .YS (\eps[12] [13]));
  FAX1 \genblk1[12].inst_SUB_UNS_OP_g1559 (.A (\eps[11] [12]), .B
       (\genblk1[12].inst_SUB_UNS_OP_n_858 ), .C
       (\genblk1[12].inst_SUB_UNS_OP_n_839 ), .YC
       (\genblk1[12].inst_SUB_UNS_OP_n_837 ), .YS (\eps[12] [12]));
  FAX1 \genblk1[12].inst_SUB_UNS_OP_g1560 (.A (\eps[11] [11]), .B
       (\genblk1[12].inst_SUB_UNS_OP_n_876 ), .C
       (\genblk1[12].inst_SUB_UNS_OP_n_841 ), .YC
       (\genblk1[12].inst_SUB_UNS_OP_n_839 ), .YS (\eps[12] [11]));
  FAX1 \genblk1[12].inst_SUB_UNS_OP_g1561 (.A (\eps[11] [10]), .B
       (\genblk1[12].inst_SUB_UNS_OP_n_867 ), .C
       (\genblk1[12].inst_SUB_UNS_OP_n_843 ), .YC
       (\genblk1[12].inst_SUB_UNS_OP_n_841 ), .YS (\eps[12] [10]));
  INVX1 \genblk1[12].inst_SUB_UNS_OP_g1562 (.A
       (\genblk1[12].inst_SUB_UNS_OP_n_844 ), .Y (\eps[12] [9]));
  INVX1 \genblk1[12].inst_SUB_UNS_OP_g1563 (.A
       (\genblk1[12].inst_SUB_UNS_OP_n_845 ), .Y
       (\genblk1[12].inst_SUB_UNS_OP_n_843 ));
  HAX1 \genblk1[12].inst_SUB_UNS_OP_g1564 (.A
       (\genblk1[12].inst_SUB_UNS_OP_n_854 ), .B
       (\genblk1[12].inst_SUB_UNS_OP_n_848 ), .YC
       (\genblk1[12].inst_SUB_UNS_OP_n_845 ), .YS
       (\genblk1[12].inst_SUB_UNS_OP_n_844 ));
  INVX1 \genblk1[12].inst_SUB_UNS_OP_g1565 (.A
       (\genblk1[12].inst_SUB_UNS_OP_n_847 ), .Y (\eps[12] [8]));
  HAX1 \genblk1[12].inst_SUB_UNS_OP_g1566 (.A
       (\genblk1[12].inst_SUB_UNS_OP_n_865 ), .B (result[4]), .YC
       (\genblk1[12].inst_SUB_UNS_OP_n_848 ), .YS
       (\genblk1[12].inst_SUB_UNS_OP_n_847 ));
  OR2X1 \genblk1[12].inst_SUB_UNS_OP_g1567 (.A
       (\genblk1[12].inst_SUB_UNS_OP_n_850 ), .B
       (\genblk1[12].inst_SUB_UNS_OP_n_852 ), .Y
       (\genblk1[12].inst_SUB_UNS_OP_n_849 ));
  AND2X1 \genblk1[12].inst_SUB_UNS_OP_g1568 (.A
       (\genblk1[12].inst_SUB_UNS_OP_n_871 ), .B (\eps[11] [20]), .Y
       (\genblk1[12].inst_SUB_UNS_OP_n_850 ));
  AND2X1 \genblk1[12].inst_SUB_UNS_OP_g1570 (.A
       (\genblk1[12].inst_n_709 ), .B
       (\genblk1[12].inst_SUB_UNS_OP_n_869 ), .Y
       (\genblk1[12].inst_SUB_UNS_OP_n_852 ));
  INVX1 \genblk1[12].inst_SUB_UNS_OP_g1571 (.A (\genblk1[12].inst_n_710
       ), .Y (\genblk1[12].inst_SUB_UNS_OP_n_853 ));
  INVX1 \genblk1[12].inst_SUB_UNS_OP_g1572 (.A (query[9]), .Y
       (\genblk1[12].inst_SUB_UNS_OP_n_854 ));
  INVX1 \genblk1[12].inst_SUB_UNS_OP_g1574 (.A (\genblk1[12].inst_n_713
       ), .Y (\genblk1[12].inst_SUB_UNS_OP_n_857 ));
  INVX1 \genblk1[12].inst_SUB_UNS_OP_g1575 (.A (\genblk1[12].inst_n_717
       ), .Y (\genblk1[12].inst_SUB_UNS_OP_n_858 ));
  INVX1 \genblk1[12].inst_SUB_UNS_OP_g1576 (.A (\genblk1[12].inst_n_711
       ), .Y (\genblk1[12].inst_SUB_UNS_OP_n_859 ));
  INVX1 \genblk1[12].inst_SUB_UNS_OP_g1578 (.A (\genblk1[12].inst_n_712
       ), .Y (\genblk1[12].inst_SUB_UNS_OP_n_862 ));
  INVX1 \genblk1[12].inst_SUB_UNS_OP_g1580 (.A (query[8]), .Y
       (\genblk1[12].inst_SUB_UNS_OP_n_865 ));
  INVX1 \genblk1[12].inst_SUB_UNS_OP_g1581 (.A (\genblk1[12].inst_n_714
       ), .Y (\genblk1[12].inst_SUB_UNS_OP_n_866 ));
  INVX1 \genblk1[12].inst_SUB_UNS_OP_g1582 (.A (\genblk1[12].inst_n_719
       ), .Y (\genblk1[12].inst_SUB_UNS_OP_n_867 ));
  INVX1 \genblk1[12].inst_SUB_UNS_OP_g1583 (.A (\eps[11] [20]), .Y
       (\genblk1[12].inst_SUB_UNS_OP_n_869 ));
  INVX1 \genblk1[12].inst_SUB_UNS_OP_g1584 (.A (\genblk1[12].inst_n_709
       ), .Y (\genblk1[12].inst_SUB_UNS_OP_n_871 ));
  INVX1 \genblk1[12].inst_SUB_UNS_OP_g1585 (.A (\genblk1[12].inst_n_716
       ), .Y (\genblk1[12].inst_SUB_UNS_OP_n_873 ));
  INVX1 \genblk1[12].inst_SUB_UNS_OP_g1586 (.A (\genblk1[12].inst_n_715
       ), .Y (\genblk1[12].inst_SUB_UNS_OP_n_874 ));
  INVX1 \genblk1[12].inst_SUB_UNS_OP_g1587 (.A (\genblk1[12].inst_n_718
       ), .Y (\genblk1[12].inst_SUB_UNS_OP_n_876 ));
  OR2X1 \genblk1[11].inst_SUB_UNS_OP_g1377 (.A (1'b0), .B (1'b0), .Y
       (\eps[11] [31]));
  FAX1 \genblk1[11].inst_SUB_UNS_OP_g1384 (.A (\eps[10] [21]), .B
       (\genblk1[11].inst_SUB_UNS_OP_n_800 ), .C
       (\genblk1[11].inst_SUB_UNS_OP_n_774 ), .YC
       (\genblk1[11].inst_SUB_UNS_OP_n_771 ), .YS (\eps[11] [21]));
  FAX1 \genblk1[11].inst_SUB_UNS_OP_g1385 (.A (\eps[10] [20]), .B
       (\genblk1[11].inst_SUB_UNS_OP_n_811 ), .C
       (\genblk1[11].inst_SUB_UNS_OP_n_776 ), .YC
       (\genblk1[11].inst_SUB_UNS_OP_n_774 ), .YS (\eps[11] [20]));
  FAX1 \genblk1[11].inst_SUB_UNS_OP_g1386 (.A (\eps[10] [19]), .B
       (\genblk1[11].inst_SUB_UNS_OP_n_810 ), .C
       (\genblk1[11].inst_SUB_UNS_OP_n_778 ), .YC
       (\genblk1[11].inst_SUB_UNS_OP_n_776 ), .YS (\eps[11] [19]));
  FAX1 \genblk1[11].inst_SUB_UNS_OP_g1387 (.A (\eps[10] [18]), .B
       (\genblk1[11].inst_SUB_UNS_OP_n_798 ), .C
       (\genblk1[11].inst_SUB_UNS_OP_n_780 ), .YC
       (\genblk1[11].inst_SUB_UNS_OP_n_778 ), .YS (\eps[11] [18]));
  FAX1 \genblk1[11].inst_SUB_UNS_OP_g1388 (.A (\eps[10] [17]), .B
       (\genblk1[11].inst_SUB_UNS_OP_n_808 ), .C
       (\genblk1[11].inst_SUB_UNS_OP_n_782 ), .YC
       (\genblk1[11].inst_SUB_UNS_OP_n_780 ), .YS (\eps[11] [17]));
  FAX1 \genblk1[11].inst_SUB_UNS_OP_g1389 (.A (\eps[10] [16]), .B
       (\genblk1[11].inst_SUB_UNS_OP_n_804 ), .C
       (\genblk1[11].inst_SUB_UNS_OP_n_784 ), .YC
       (\genblk1[11].inst_SUB_UNS_OP_n_782 ), .YS (\eps[11] [16]));
  FAX1 \genblk1[11].inst_SUB_UNS_OP_g1390 (.A (\eps[10] [15]), .B
       (\genblk1[11].inst_SUB_UNS_OP_n_803 ), .C
       (\genblk1[11].inst_SUB_UNS_OP_n_786 ), .YC
       (\genblk1[11].inst_SUB_UNS_OP_n_784 ), .YS (\eps[11] [15]));
  FAX1 \genblk1[11].inst_SUB_UNS_OP_g1391 (.A (\eps[10] [14]), .B
       (\genblk1[11].inst_SUB_UNS_OP_n_806 ), .C
       (\genblk1[11].inst_SUB_UNS_OP_n_788 ), .YC
       (\genblk1[11].inst_SUB_UNS_OP_n_786 ), .YS (\eps[11] [14]));
  FAX1 \genblk1[11].inst_SUB_UNS_OP_g1392 (.A (\eps[10] [13]), .B
       (\genblk1[11].inst_SUB_UNS_OP_n_805 ), .C
       (\genblk1[11].inst_SUB_UNS_OP_n_790 ), .YC
       (\genblk1[11].inst_SUB_UNS_OP_n_788 ), .YS (\eps[11] [13]));
  FAX1 \genblk1[11].inst_SUB_UNS_OP_g1393 (.A (\eps[10] [12]), .B
       (\genblk1[11].inst_SUB_UNS_OP_n_802 ), .C
       (\genblk1[11].inst_SUB_UNS_OP_n_792 ), .YC
       (\genblk1[11].inst_SUB_UNS_OP_n_790 ), .YS (\eps[11] [12]));
  INVX1 \genblk1[11].inst_SUB_UNS_OP_g1394 (.A
       (\genblk1[11].inst_SUB_UNS_OP_n_793 ), .Y (\eps[11] [11]));
  INVX1 \genblk1[11].inst_SUB_UNS_OP_g1395 (.A
       (\genblk1[11].inst_SUB_UNS_OP_n_794 ), .Y
       (\genblk1[11].inst_SUB_UNS_OP_n_792 ));
  HAX1 \genblk1[11].inst_SUB_UNS_OP_g1396 (.A
       (\genblk1[11].inst_SUB_UNS_OP_n_807 ), .B
       (\genblk1[11].inst_SUB_UNS_OP_n_797 ), .YC
       (\genblk1[11].inst_SUB_UNS_OP_n_794 ), .YS
       (\genblk1[11].inst_SUB_UNS_OP_n_793 ));
  INVX1 \genblk1[11].inst_SUB_UNS_OP_g1397 (.A
       (\genblk1[11].inst_SUB_UNS_OP_n_796 ), .Y (\eps[11] [10]));
  HAX1 \genblk1[11].inst_SUB_UNS_OP_g1398 (.A
       (\genblk1[11].inst_SUB_UNS_OP_n_801 ), .B (result[5]), .YC
       (\genblk1[11].inst_SUB_UNS_OP_n_797 ), .YS
       (\genblk1[11].inst_SUB_UNS_OP_n_796 ));
  INVX1 \genblk1[11].inst_SUB_UNS_OP_g1399 (.A (\genblk1[11].inst_n_711
       ), .Y (\genblk1[11].inst_SUB_UNS_OP_n_798 ));
  INVX1 \genblk1[11].inst_SUB_UNS_OP_g1400 (.A (\genblk1[11].inst_n_708
       ), .Y (\genblk1[11].inst_SUB_UNS_OP_n_800 ));
  INVX1 \genblk1[11].inst_SUB_UNS_OP_g1401 (.A (query[10]), .Y
       (\genblk1[11].inst_SUB_UNS_OP_n_801 ));
  INVX1 \genblk1[11].inst_SUB_UNS_OP_g1402 (.A (\genblk1[11].inst_n_717
       ), .Y (\genblk1[11].inst_SUB_UNS_OP_n_802 ));
  INVX1 \genblk1[11].inst_SUB_UNS_OP_g1403 (.A (\genblk1[11].inst_n_714
       ), .Y (\genblk1[11].inst_SUB_UNS_OP_n_803 ));
  INVX1 \genblk1[11].inst_SUB_UNS_OP_g1404 (.A (\genblk1[11].inst_n_713
       ), .Y (\genblk1[11].inst_SUB_UNS_OP_n_804 ));
  INVX1 \genblk1[11].inst_SUB_UNS_OP_g1405 (.A (\genblk1[11].inst_n_716
       ), .Y (\genblk1[11].inst_SUB_UNS_OP_n_805 ));
  INVX1 \genblk1[11].inst_SUB_UNS_OP_g1406 (.A (\genblk1[11].inst_n_715
       ), .Y (\genblk1[11].inst_SUB_UNS_OP_n_806 ));
  INVX1 \genblk1[11].inst_SUB_UNS_OP_g1407 (.A (query[11]), .Y
       (\genblk1[11].inst_SUB_UNS_OP_n_807 ));
  INVX1 \genblk1[11].inst_SUB_UNS_OP_g1408 (.A (\genblk1[11].inst_n_712
       ), .Y (\genblk1[11].inst_SUB_UNS_OP_n_808 ));
  INVX1 \genblk1[11].inst_SUB_UNS_OP_g1409 (.A (\genblk1[11].inst_n_710
       ), .Y (\genblk1[11].inst_SUB_UNS_OP_n_810 ));
  INVX1 \genblk1[11].inst_SUB_UNS_OP_g1410 (.A (\genblk1[11].inst_n_709
       ), .Y (\genblk1[11].inst_SUB_UNS_OP_n_811 ));
  FAX1 \genblk1[10].inst_SUB_UNS_OP_g1246 (.A (\eps[9] [22]), .B
       (\genblk1[10].inst_SUB_UNS_OP_n_760 ), .C
       (\genblk1[10].inst_SUB_UNS_OP_n_738 ), .YC
       (\genblk1[10].inst_SUB_UNS_OP_n_736 ), .YS (\eps[10] [22]));
  FAX1 \genblk1[10].inst_SUB_UNS_OP_g1247 (.A (\eps[9] [21]), .B
       (\genblk1[10].inst_SUB_UNS_OP_n_763 ), .C
       (\genblk1[10].inst_SUB_UNS_OP_n_740 ), .YC
       (\genblk1[10].inst_SUB_UNS_OP_n_738 ), .YS (\eps[10] [21]));
  FAX1 \genblk1[10].inst_SUB_UNS_OP_g1248 (.A (\eps[9] [20]), .B
       (\genblk1[10].inst_SUB_UNS_OP_n_771 ), .C
       (\genblk1[10].inst_SUB_UNS_OP_n_742 ), .YC
       (\genblk1[10].inst_SUB_UNS_OP_n_740 ), .YS (\eps[10] [20]));
  FAX1 \genblk1[10].inst_SUB_UNS_OP_g1249 (.A (\eps[9] [19]), .B
       (\genblk1[10].inst_SUB_UNS_OP_n_769 ), .C
       (\genblk1[10].inst_SUB_UNS_OP_n_744 ), .YC
       (\genblk1[10].inst_SUB_UNS_OP_n_742 ), .YS (\eps[10] [19]));
  FAX1 \genblk1[10].inst_SUB_UNS_OP_g1250 (.A (\eps[9] [18]), .B
       (\genblk1[10].inst_SUB_UNS_OP_n_768 ), .C
       (\genblk1[10].inst_SUB_UNS_OP_n_746 ), .YC
       (\genblk1[10].inst_SUB_UNS_OP_n_744 ), .YS (\eps[10] [18]));
  FAX1 \genblk1[10].inst_SUB_UNS_OP_g1251 (.A (\eps[9] [17]), .B
       (\genblk1[10].inst_SUB_UNS_OP_n_767 ), .C
       (\genblk1[10].inst_SUB_UNS_OP_n_748 ), .YC
       (\genblk1[10].inst_SUB_UNS_OP_n_746 ), .YS (\eps[10] [17]));
  FAX1 \genblk1[10].inst_SUB_UNS_OP_g1252 (.A (\eps[9] [16]), .B
       (\genblk1[10].inst_SUB_UNS_OP_n_765 ), .C
       (\genblk1[10].inst_SUB_UNS_OP_n_750 ), .YC
       (\genblk1[10].inst_SUB_UNS_OP_n_748 ), .YS (\eps[10] [16]));
  FAX1 \genblk1[10].inst_SUB_UNS_OP_g1253 (.A (\eps[9] [15]), .B
       (\genblk1[10].inst_SUB_UNS_OP_n_766 ), .C
       (\genblk1[10].inst_SUB_UNS_OP_n_752 ), .YC
       (\genblk1[10].inst_SUB_UNS_OP_n_750 ), .YS (\eps[10] [15]));
  FAX1 \genblk1[10].inst_SUB_UNS_OP_g1254 (.A (\eps[9] [14]), .B
       (\genblk1[10].inst_SUB_UNS_OP_n_764 ), .C
       (\genblk1[10].inst_SUB_UNS_OP_n_754 ), .YC
       (\genblk1[10].inst_SUB_UNS_OP_n_752 ), .YS (\eps[10] [14]));
  INVX1 \genblk1[10].inst_SUB_UNS_OP_g1255 (.A
       (\genblk1[10].inst_SUB_UNS_OP_n_755 ), .Y (\eps[10] [13]));
  INVX1 \genblk1[10].inst_SUB_UNS_OP_g1256 (.A
       (\genblk1[10].inst_SUB_UNS_OP_n_756 ), .Y
       (\genblk1[10].inst_SUB_UNS_OP_n_754 ));
  HAX1 \genblk1[10].inst_SUB_UNS_OP_g1257 (.A
       (\genblk1[10].inst_SUB_UNS_OP_n_770 ), .B
       (\genblk1[10].inst_SUB_UNS_OP_n_759 ), .YC
       (\genblk1[10].inst_SUB_UNS_OP_n_756 ), .YS
       (\genblk1[10].inst_SUB_UNS_OP_n_755 ));
  INVX1 \genblk1[10].inst_SUB_UNS_OP_g1258 (.A
       (\genblk1[10].inst_SUB_UNS_OP_n_758 ), .Y (\eps[10] [12]));
  HAX1 \genblk1[10].inst_SUB_UNS_OP_g1259 (.A
       (\genblk1[10].inst_SUB_UNS_OP_n_761 ), .B (result[6]), .YC
       (\genblk1[10].inst_SUB_UNS_OP_n_759 ), .YS
       (\genblk1[10].inst_SUB_UNS_OP_n_758 ));
  INVX1 \genblk1[10].inst_SUB_UNS_OP_g1260 (.A (\genblk1[10].inst_n_707
       ), .Y (\genblk1[10].inst_SUB_UNS_OP_n_760 ));
  INVX1 \genblk1[10].inst_SUB_UNS_OP_g1261 (.A (query[12]), .Y
       (\genblk1[10].inst_SUB_UNS_OP_n_761 ));
  INVX1 \genblk1[10].inst_SUB_UNS_OP_g1263 (.A (\genblk1[10].inst_n_708
       ), .Y (\genblk1[10].inst_SUB_UNS_OP_n_763 ));
  INVX1 \genblk1[10].inst_SUB_UNS_OP_g1264 (.A (\genblk1[10].inst_n_715
       ), .Y (\genblk1[10].inst_SUB_UNS_OP_n_764 ));
  INVX1 \genblk1[10].inst_SUB_UNS_OP_g1265 (.A (\genblk1[10].inst_n_713
       ), .Y (\genblk1[10].inst_SUB_UNS_OP_n_765 ));
  INVX1 \genblk1[10].inst_SUB_UNS_OP_g1266 (.A (\genblk1[10].inst_n_714
       ), .Y (\genblk1[10].inst_SUB_UNS_OP_n_766 ));
  INVX1 \genblk1[10].inst_SUB_UNS_OP_g1267 (.A (\genblk1[10].inst_n_712
       ), .Y (\genblk1[10].inst_SUB_UNS_OP_n_767 ));
  INVX1 \genblk1[10].inst_SUB_UNS_OP_g1268 (.A (\genblk1[10].inst_n_711
       ), .Y (\genblk1[10].inst_SUB_UNS_OP_n_768 ));
  INVX1 \genblk1[10].inst_SUB_UNS_OP_g1269 (.A (\genblk1[10].inst_n_710
       ), .Y (\genblk1[10].inst_SUB_UNS_OP_n_769 ));
  INVX1 \genblk1[10].inst_SUB_UNS_OP_g1270 (.A (query[13]), .Y
       (\genblk1[10].inst_SUB_UNS_OP_n_770 ));
  INVX1 \genblk1[10].inst_SUB_UNS_OP_g1271 (.A (\genblk1[10].inst_n_709
       ), .Y (\genblk1[10].inst_SUB_UNS_OP_n_771 ));
endmodule

